
module MUX21_GENERIC_N4_42 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_168 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_167 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_166 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_165 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n2) );
endmodule


module MUX21_GENERIC_N4_17 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_68 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_67 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_66 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_65 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n2) );
endmodule


module MUX21_GENERIC_N4_15 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_60 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_59 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_58 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_57 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_12 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_48 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_47 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_46 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_45 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_11 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_44 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_43 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_42 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_41 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_62 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_248 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_247 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_246 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_245 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_61 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_244 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_243 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_242 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_241 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_60 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_240 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_239 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_238 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_237 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_59 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_236 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_235 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_234 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_233 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_58 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_232 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_231 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_230 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_229 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_57 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_228 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_227 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_226 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_225 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_50 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_200 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_199 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_198 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_197 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_49 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_196 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_195 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_194 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_193 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_41 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_164 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_163 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_162 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_161 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_33 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_132 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_131 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_130 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_129 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_24 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_96 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_95 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_94 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_93 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_16 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_64 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_63 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_62 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_61 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_8 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_32 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_31 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_30 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_29 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_7 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_28 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_27 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_26 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_25 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_12 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_11 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_10 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_9 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_8 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_7 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_6 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_5 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_64 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_256 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_255 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_254 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_253 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_48 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_192 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_191 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_190 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_189 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_47 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_188 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_187 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_186 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_185 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_96 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_95 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSAdd_N4_49 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_98 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_97 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_49 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_8 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_16 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_15 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_8 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genP_198 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  NAND2_X1 U2 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U3 ( .A(G1), .ZN(n8) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_193 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  NAND2_X1 U2 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U3 ( .A(G1), .ZN(n8) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_171 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_144 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  INV_X1 U1 ( .A(G1), .ZN(n8) );
  AND2_X1 U2 ( .A1(P0), .A2(P1), .ZN(Pout) );
  NAND2_X1 U3 ( .A1(n8), .A2(n7), .ZN(Gout) );
  NAND2_X1 U4 ( .A1(G0), .A2(P1), .ZN(n7) );
endmodule


module genP_85 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(n8), .A2(n7), .ZN(Gout) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_156 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_131 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_98 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_72 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_63 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_58 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net225014, net232817, n6;
  assign Pout = net232817;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net232817) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(net225014) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(net225014), .ZN(Gout) );
endmodule


module genP_213 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_212 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_211 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_209 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_208 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_207 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_204 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_202 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_201 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_199 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_197 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_196 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_194 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_191 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_190 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_186 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_181 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_180 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_179 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_178 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_177 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_170 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_169 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_159 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_158 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_154 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_153 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_151 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_150 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_143 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_142 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_137 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_133 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_132 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_129 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net226160, net232816, n6;
  assign Pout = net232816;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net232816) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(net226160) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(net226160), .ZN(Gout) );
endmodule


module genP_128 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_126 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_124 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_123 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_115 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_105 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_104 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_103 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_97 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_83 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_81 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_74 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_61 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_59 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_51 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_50 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_49 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_47 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_46 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_27 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_210 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_206 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_205 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_203 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_195 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_192 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_166 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_164 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_161 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_155 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_152 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(n6), .A2(G1), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_110 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_107 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_80 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_54 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_53 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_26 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_24 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genP_75 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_21 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_183 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_174 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_130 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_127 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_108 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_102 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_101 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_100 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_73 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_71 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net225048, net238615, n6;
  assign Pout = net238615;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net238615) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(net225048) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(net225048), .A2(n6), .ZN(Gout) );
endmodule


module genP_45 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_42 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_25 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_22 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_18 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_17 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_16 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_15 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X2 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_175 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_165 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_149 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_148 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_138 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_122 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_121 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_111 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_95 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_94 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_84 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_68 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_67 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_41 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_40 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_14 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_13 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_134 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_10 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_117 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  NAND2_X1 U2 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U3 ( .A(G1), .ZN(n8) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_62 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net225025, net233213, n6;
  assign Pout = net233213;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net233213) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(net225025) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(net225025), .ZN(Gout) );
endmodule


module genP_35 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_34 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net180042, net232910, net224494, n6;
  assign Gout = net180042;
  assign Pout = net232910;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net232910) );
  NAND2_X1 U2 ( .A1(G0), .A2(P1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(net224494), .ZN(net180042) );
  INV_X1 U4 ( .A(G1), .ZN(net224494) );
endmodule


module genP_8 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(G0), .A2(P1), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_36 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  NAND2_X1 U1 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  AND2_X1 U4 ( .A1(P0), .A2(P1), .ZN(Pout) );
endmodule


module genP_31 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(n8), .A2(n7), .ZN(Gout) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_11 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  NAND2_X1 U2 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U3 ( .A(G1), .ZN(n8) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_4 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(n8), .A2(n7), .ZN(Gout) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_141 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_114 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_109 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_87 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_82 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_60 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_57 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_33 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_30 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_28 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_6 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_3 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_167 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_162 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_160 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_147 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_146 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(G0), .A2(P1), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_140 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_135 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_125 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_119 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_118 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net226131, net232815, n6;
  assign Pout = net232815;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net232815) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(net226131) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(net226131), .A2(n6), .ZN(Gout) );
endmodule


module genP_116 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_113 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net226117, net239227, n6;
  assign Pout = net239227;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(net239227) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(net226117) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(net226117), .ZN(Gout) );
endmodule


module genP_106 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_96 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_93 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_91 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_89 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_88 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  OR2_X2 U1 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_86 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_79 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_78 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_77 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_70 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_69 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_66 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_56 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  OR2_X1 U1 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n6) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_52 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_48 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_44 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_39 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_37 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(G0), .A2(P1), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_32 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_29 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net180021, net241284, n6, n7;
  assign Gout = net180021;
  assign Pout = net241284;

  NAND2_X1 U1 ( .A1(n6), .A2(n7), .ZN(net180021) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n7) );
  INV_X1 U3 ( .A(G1), .ZN(n6) );
  AND2_X1 U4 ( .A1(P0), .A2(P1), .ZN(net241284) );
endmodule


module genP_23 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_19 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_12 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_7 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X2 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_5 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_2 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_136 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_55 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_1 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genG_70 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  INV_X1 U1 ( .A(G1), .ZN(n6) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_68 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  INV_X1 U1 ( .A(G1), .ZN(n6) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_65 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  INV_X1 U1 ( .A(G1), .ZN(n6) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_54 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_51 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net182392, n4, n5;
  assign Gout = net182392;

  NAND2_X2 U1 ( .A1(n5), .A2(n4), .ZN(net182392) );
  INV_X1 U2 ( .A(G1), .ZN(n4) );
  NAND2_X1 U3 ( .A1(G0), .A2(P1), .ZN(n5) );
endmodule


module genG_67 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_66 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_64 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_57 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_56 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_47 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_38 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_22 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X2 U1 ( .A1(n5), .A2(n6), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n5) );
endmodule


module genG_36 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_27 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_18 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_9 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genG_53 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4, n5;

  NAND2_X2 U1 ( .A1(n5), .A2(n4), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_50 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net182389, n4;
  assign Gout = net182389;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(net182389) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_44 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4, n5;

  INV_X1 U1 ( .A(G1), .ZN(n5) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
  NAND2_X2 U3 ( .A1(n5), .A2(n4), .ZN(Gout) );
endmodule


module genG_43 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4, n5;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_33 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(G0), .A2(P1), .ZN(n4) );
endmodule


module genG_30 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_29 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_24 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_21 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net180606, n4;
  assign Gout = net180606;

  AND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n4) );
  OR2_X2 U2 ( .A1(n4), .A2(G1), .ZN(net180606) );
endmodule


module genG_20 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_16 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_7 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_3 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_48 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_41 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net181798, n4;
  assign Gout = net181798;

  AND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n4) );
  OR2_X2 U2 ( .A1(G1), .A2(n4), .ZN(net181798) );
endmodule


module genG_39 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4, n5;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n5) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_34 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_32 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net181207, n4;
  assign Gout = net181207;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(net181207) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_26 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4, n5;

  INV_X1 U1 ( .A(G1), .ZN(n5) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
  NAND2_X2 U3 ( .A1(n5), .A2(n4), .ZN(Gout) );
endmodule


module genG_25 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_23 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_17 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4, n5;

  INV_X1 U1 ( .A(G1), .ZN(n5) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
  NAND2_X2 U3 ( .A1(n5), .A2(n4), .ZN(Gout) );
endmodule


module genG_15 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_14 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_12 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_11 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net180012, n4;
  assign Gout = net180012;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(net180012) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_5 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_2 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net179421, n4;
  assign Gout = net179421;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(net179421) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_46 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n4) );
endmodule


module genG_37 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n4) );
endmodule


module genG_28 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n4) );
endmodule


module genG_19 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n4) );
endmodule


module genG_10 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n4) );
endmodule


module genG_1 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n4) );
endmodule


module PGblock_209 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_208 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_206 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(b), .ZN(n3) );
  XNOR2_X1 U3 ( .A(a), .B(n3), .ZN(p) );
endmodule


module PGblock_201 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_199 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_198 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_197 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_196 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_195 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_194 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_193 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_192 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_191 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_180 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n5;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n5) );
  XNOR2_X1 U3 ( .A(b), .B(n5), .ZN(p) );
endmodule


module PGblock_143 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_108 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_164 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_140 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_109 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_104 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  CLKBUF_X1 U1 ( .A(b), .Z(n2) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U3 ( .A1(n2), .A2(a), .ZN(g) );
endmodule


module PGblock_98 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_236 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_234 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_232 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_224 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_220 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_217 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_212 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_178 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_177 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_174 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_171 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_170 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_169 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_162 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_155 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_147 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_131 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_124 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_116 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_112 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_100 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_93 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_85 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_77 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_69 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_68 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_46 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_31 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_30 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_23 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_19 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_15 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_25 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_21 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_13 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_246 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_245 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_244 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_243 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_242 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_241 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_239 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_238 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_237 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_235 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_233 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_231 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_230 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_229 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_228 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_227 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_226 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_225 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_223 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_222 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_221 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_219 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_218 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_214 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_205 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  CLKBUF_X1 U1 ( .A(b), .Z(n2) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U3 ( .A1(a), .A2(n2), .ZN(g) );
endmodule


module PGblock_204 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_203 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_183 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_182 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_179 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_168 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_167 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_166 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_165 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_163 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_161 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_160 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_152 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_151 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_148 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_146 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_142 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_138 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_135 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_134 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_132 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_130 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_129 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_121 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_120 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_117 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_101 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_99 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_90 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_86 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_82 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_80 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_78 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_76 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_61 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_55 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_51 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_47 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_45 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_44 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_37 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_28 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_27 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_26 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_24 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_22 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_20 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_18 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_14 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_10 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n2;

  INV_X1 U1 ( .A(a), .ZN(n2) );
  XNOR2_X1 U2 ( .A(b), .B(n2), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_141 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   net238672, n3;
  assign g = net238672;

  XNOR2_X1 U1 ( .A(b), .B(n3), .ZN(p) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(net238672) );
endmodule


module PGblock_133 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_72 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_42 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_41 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_11 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_9 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  AND2_X1 U3 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_181 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_154 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_153 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_149 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_144 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_123 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_119 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_118 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_115 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_113 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_111 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_107 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_105 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_92 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_91 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_89 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_88 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_84 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_81 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_70 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_62 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_60 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_59 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_58 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_57 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_54 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_53 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_52 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_50 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_49 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_48 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_43 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_39 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_17 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4, n5;

  AND2_X1 U1 ( .A1(a), .A2(n4), .ZN(g) );
  CLKBUF_X1 U2 ( .A(b), .Z(n4) );
  INV_X1 U3 ( .A(a), .ZN(n5) );
  XNOR2_X1 U4 ( .A(b), .B(n5), .ZN(p) );
endmodule


module PGblock_12 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_8 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_150 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_139 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_136 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_122 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_114 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_110 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   net239234, n3;
  assign g = net239234;

  XNOR2_X1 U1 ( .A(b), .B(n3), .ZN(p) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(net239234) );
endmodule


module PGblock_106 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_83 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_74 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_56 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_38 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   net239229, n3;
  assign g = net239229;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(net239229) );
endmodule


module PGblock_7 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_102 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  INV_X1 U1 ( .A(a), .ZN(n4) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_75 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_73 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_67 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4, n5;

  INV_X1 U1 ( .A(a), .ZN(n5) );
  AND2_X1 U2 ( .A1(n4), .A2(a), .ZN(g) );
  CLKBUF_X1 U3 ( .A(b), .Z(n4) );
  XNOR2_X1 U4 ( .A(b), .B(n5), .ZN(p) );
endmodule


module PGblock_40 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  CLKBUF_X1 U1 ( .A(b), .Z(n3) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U3 ( .A1(n3), .A2(a), .ZN(g) );
endmodule


module PGblock_36 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_6 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_5 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   net239221, n3, n4;
  assign g = net239221;

  INV_X1 U1 ( .A(a), .ZN(n3) );
  XNOR2_X1 U2 ( .A(b), .B(n3), .ZN(p) );
  CLKBUF_X1 U3 ( .A(b), .Z(n4) );
  AND2_X1 U4 ( .A1(n4), .A2(a), .ZN(net239221) );
endmodule


module PGblock_189 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_188 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_187 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_159 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_158 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_157 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_156 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_128 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_127 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_126 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_125 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_97 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_96 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_95 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_94 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_66 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_65 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_64 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_63 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_35 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_34 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_33 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_32 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module Gstart_5 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module Gstart_4 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module Gstart_3 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module Gstart_2 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module Gstart_1 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module Boothencoder_4 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   n9, n10, n11;

  OAI21_X1 U1 ( .B1(B[0]), .B2(B[1]), .A(n11), .ZN(n10) );
  NAND2_X1 U2 ( .A1(B[1]), .A2(B[0]), .ZN(n11) );
  AND3_X1 U3 ( .A1(n11), .A2(B[2]), .A3(n10), .ZN(S[2]) );
  AOI21_X1 U4 ( .B1(n11), .B2(n10), .A(B[2]), .ZN(S[0]) );
  MUX2_X1 U5 ( .A(n11), .B(n10), .S(B[2]), .Z(n9) );
  INV_X1 U6 ( .A(n9), .ZN(S[1]) );
endmodule


module Boothencoder_3 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   n9, n10, n11;

  OAI21_X1 U1 ( .B1(B[0]), .B2(B[1]), .A(n11), .ZN(n10) );
  NAND2_X1 U2 ( .A1(B[1]), .A2(B[0]), .ZN(n11) );
  AND3_X1 U3 ( .A1(n11), .A2(B[2]), .A3(n10), .ZN(S[2]) );
  AOI21_X1 U4 ( .B1(n11), .B2(n10), .A(B[2]), .ZN(S[0]) );
  MUX2_X1 U5 ( .A(n11), .B(n10), .S(B[2]), .Z(n9) );
  INV_X1 U6 ( .A(n9), .ZN(S[1]) );
endmodule


module Boothencoder_2 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   n9, n10, n11;

  OAI21_X1 U1 ( .B1(B[0]), .B2(B[1]), .A(n11), .ZN(n10) );
  NAND2_X1 U2 ( .A1(B[1]), .A2(B[0]), .ZN(n11) );
  AND3_X1 U3 ( .A1(n11), .A2(B[2]), .A3(n10), .ZN(S[2]) );
  AOI21_X1 U4 ( .B1(n11), .B2(n10), .A(B[2]), .ZN(S[0]) );
  MUX2_X1 U5 ( .A(n11), .B(n10), .S(B[2]), .Z(n9) );
  INV_X1 U6 ( .A(n9), .ZN(S[1]) );
endmodule


module Boothencoder_1 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   n9, n10, n11;

  OAI21_X1 U1 ( .B1(B[0]), .B2(B[1]), .A(n11), .ZN(n10) );
  NAND2_X1 U2 ( .A1(B[1]), .A2(B[0]), .ZN(n11) );
  AND3_X1 U3 ( .A1(n11), .A2(B[2]), .A3(n10), .ZN(S[2]) );
  AOI21_X1 U4 ( .B1(n11), .B2(n10), .A(B[2]), .ZN(S[0]) );
  MUX2_X1 U5 ( .A(n11), .B(n10), .S(B[2]), .Z(n9) );
  INV_X1 U6 ( .A(n9), .ZN(S[1]) );
endmodule


module ND2_2825 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2822 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2819 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2816 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2813 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2810 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2807 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2804 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2801 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2798 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2795 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2761 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2758 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2739 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2738 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2737 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2736 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2735 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2734 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2733 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2732 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2731 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2730 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2729 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2728 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2727 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2726 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2725 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2723 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2720 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2717 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2714 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2711 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1728 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1727 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1726 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1725 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1724 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1723 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1722 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1721 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1720 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1719 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1718 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1717 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1716 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1715 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1714 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1713 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1712 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1711 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1710 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1709 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1708 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1707 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1706 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1705 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1704 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1703 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1702 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1701 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1700 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1699 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1698 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1697 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1696 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1695 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1694 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1693 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1692 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1691 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1690 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1689 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1688 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1687 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_934 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_928 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_925 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_916 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_913 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_910 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_907 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_904 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_901 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_886 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_880 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_877 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_874 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_871 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_868 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_865 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_838 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_835 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_832 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_829 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_826 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_820 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_817 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_805 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_802 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_784 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_781 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_778 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_775 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_772 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_769 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_661 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_601 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_72 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_69 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_60 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_57 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_54 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_48 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_45 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_44 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_36 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_33 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_24 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_21 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_18 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_12 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_9 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_6 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_3 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2826 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2824 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2823 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2821 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2820 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2818 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2817 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2815 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2814 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2812 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2811 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2809 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2808 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2806 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2805 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2803 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2802 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2800 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2799 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2797 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2796 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2794 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2793 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2792 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2791 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2790 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2789 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2788 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2787 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2786 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2785 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2784 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2783 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2782 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2781 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2780 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2779 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2778 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2777 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2776 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2775 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2774 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2773 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2772 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2771 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2770 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2769 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2768 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2767 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2766 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2765 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2764 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2763 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2762 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2760 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2759 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2757 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2756 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2755 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2754 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2753 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2752 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2751 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2750 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2749 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2748 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2747 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2746 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2745 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2744 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2743 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2742 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2741 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2740 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2724 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2722 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2721 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2719 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2718 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2716 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2715 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2713 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2712 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2710 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2709 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2708 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2707 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2706 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2705 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2704 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2703 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2702 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2701 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2700 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2699 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2698 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2697 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2696 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2695 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2694 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2693 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2692 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2691 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2690 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2689 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2688 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2687 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2670 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2664 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2660 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2659 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2636 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2633 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2632 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2630 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2629 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2627 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2564 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2553 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2552 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2541 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2540 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2539 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2528 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2525 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2519 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2516 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2515 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2513 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2468 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2456 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2444 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2212 ( A, B, Y );
  input A, B;
  output Y;
  wire   n2;

  BUF_X2 U1 ( .A(n2), .Z(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module ND2_2211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2200 ( A, B, Y );
  input A, B;
  output Y;
  wire   n2;

  BUF_X4 U1 ( .A(n2), .Z(Y) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n2) );
endmodule


module ND2_2199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2099 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2098 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2097 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2096 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2095 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2094 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2093 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2092 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2091 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2090 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2089 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2088 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2087 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2086 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2085 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2084 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2083 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2082 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2081 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2080 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2079 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2078 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2077 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2076 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2075 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2074 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2073 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2072 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2071 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2070 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2069 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2068 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2067 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2066 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2065 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2064 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2063 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2062 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2061 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2060 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2059 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2058 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2057 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2056 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2055 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2054 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2053 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2052 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2051 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2050 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2049 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2048 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2047 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2046 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2045 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2044 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2043 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2042 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2041 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2040 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2039 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2038 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2037 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2036 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2035 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2034 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_2033 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2032 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2031 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2030 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2029 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2028 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2027 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2026 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2025 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2024 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2023 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2022 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2021 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2020 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2019 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2018 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2017 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2016 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2015 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2014 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2013 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2012 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2011 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2010 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2009 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2008 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2007 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2006 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2005 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2004 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2003 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2002 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2001 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2000 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1999 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1998 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1997 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1996 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1995 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1994 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1993 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1992 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1991 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1990 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1989 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1988 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1987 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1986 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1985 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1984 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1983 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1982 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1981 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1980 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1979 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1978 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1977 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1976 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1975 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1974 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1973 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1972 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1971 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1970 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1969 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1968 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1967 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1966 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1965 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1964 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1963 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1962 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1961 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1960 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1959 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1958 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1957 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1956 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1955 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1954 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1953 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1952 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1951 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1950 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1949 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1948 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1947 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1946 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1945 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1944 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1943 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1942 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1941 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1940 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1938 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1937 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1935 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1934 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1933 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1932 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1931 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1929 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1928 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1926 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1925 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1923 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1922 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1921 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1920 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1919 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1917 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1916 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1915 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1914 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1913 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1911 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1910 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1909 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1908 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1907 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1905 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1904 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1903 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1902 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1901 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1899 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1898 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1897 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1896 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1895 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1894 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1893 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1892 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1891 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1890 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1889 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1888 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1887 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1886 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1885 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1884 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1883 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1882 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1881 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1880 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1879 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1878 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1877 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1876 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1875 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1874 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1873 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1872 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1871 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1870 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1869 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1868 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1867 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1866 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1865 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1864 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1863 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1862 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1861 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1860 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1859 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1858 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1857 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1856 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1855 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1854 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1853 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1852 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1851 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1850 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1849 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1848 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1847 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1846 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1845 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1844 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1843 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1842 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1841 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1840 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1839 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1838 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1837 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1836 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1835 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1834 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1833 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1832 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1831 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1830 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1829 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1828 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1827 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1826 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1825 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1824 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1823 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1822 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1821 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1820 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1819 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1818 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1817 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1816 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1815 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1814 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1813 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1812 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1811 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1810 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1809 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1808 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1807 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1806 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1805 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1804 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1803 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1802 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1801 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1800 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1799 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1798 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1797 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1796 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1795 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1794 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1793 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1792 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1791 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1790 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1789 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1788 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1787 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1786 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1785 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1784 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1783 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1782 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1781 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1780 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1779 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1778 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1777 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1776 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1775 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1774 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1773 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1772 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1771 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1770 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1769 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1768 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1767 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1766 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1765 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1764 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1763 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1762 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1761 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1760 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1759 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1758 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1757 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1756 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1755 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1754 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1753 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1752 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1751 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1750 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1749 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1748 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1747 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1746 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1745 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1744 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1743 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1742 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1741 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1740 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1739 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1738 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1737 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1736 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1735 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1734 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1733 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1732 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1731 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1730 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1729 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1433 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1432 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1421 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1420 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1417 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1414 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1372 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1361 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1360 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1342 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1324 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1323 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1321 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1318 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1312 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1311 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1309 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1264 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1253 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1252 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1239 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1228 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1225 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1222 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1217 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1216 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1213 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1205 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1204 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1168 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1158 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1157 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1156 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1144 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1132 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1120 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1117 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1108 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1107 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1105 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1099 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1098 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1097 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1096 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1095 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1094 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1093 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1092 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1091 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1090 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1089 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1088 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1087 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1086 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1085 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1084 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1083 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1082 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1081 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1080 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1079 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1078 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1077 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1076 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1075 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1074 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1073 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1072 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1071 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1070 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1069 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1068 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1067 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1066 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1065 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1064 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1063 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1062 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1061 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1060 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1059 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1058 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1057 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1056 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1055 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1054 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1053 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1052 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1051 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1050 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1049 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1048 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1047 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1046 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1045 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1044 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1043 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1042 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1041 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1040 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1039 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1038 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1037 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1036 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1035 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1034 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1033 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1032 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1031 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1030 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1029 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1028 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1027 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1026 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1025 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1024 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1023 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1022 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1021 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1020 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1019 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1018 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1017 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1016 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1015 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1014 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1013 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1012 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1011 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1010 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1009 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1008 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1007 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1006 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1005 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1004 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1003 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1002 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1001 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1000 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_999 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_998 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_997 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_996 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_995 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_994 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_993 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_992 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_991 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_990 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_989 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_988 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_987 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_986 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_985 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_984 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_983 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_982 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_981 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_980 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_979 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_978 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_977 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_976 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_975 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_974 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_973 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_972 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_971 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_970 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_969 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_968 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_967 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_966 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_965 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_964 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_963 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_962 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_961 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_960 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_959 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_958 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_957 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_956 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_955 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_954 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_953 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_952 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_951 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_950 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_949 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_948 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_947 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_946 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_945 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_944 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_943 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_942 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_941 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_940 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_939 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_938 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_937 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_936 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_935 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_933 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_932 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_931 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_930 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_929 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_927 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_926 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_924 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_923 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_922 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_921 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_920 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_919 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_918 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_917 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_915 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_914 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_912 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_911 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_909 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_908 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_906 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_905 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_903 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_902 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_900 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_899 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_898 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_897 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_896 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_895 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_894 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_893 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_892 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_891 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_890 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_889 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_888 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_887 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_885 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_884 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_883 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_882 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_881 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_879 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_878 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_876 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_875 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_873 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_872 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_870 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_869 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_867 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_866 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_864 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_863 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_862 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_861 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_860 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_859 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_858 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_857 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_856 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_855 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_854 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_853 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_852 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_851 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_850 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_849 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_848 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_847 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_846 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_845 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_844 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_843 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_842 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_841 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_840 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_839 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_837 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_836 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_834 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_833 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_831 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_830 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_828 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_827 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_825 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_824 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_823 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_822 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_821 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_819 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_818 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_816 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_815 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_814 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_813 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_812 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_811 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_810 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_809 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_808 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_807 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_806 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_804 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_803 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_801 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_800 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_799 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_798 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_797 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_796 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_795 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_794 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_793 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_792 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_791 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_790 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_789 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_788 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_787 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_786 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_785 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_783 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_782 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_780 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_779 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_777 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_776 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_774 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_773 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_771 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_770 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_768 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_767 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_766 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_765 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_764 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_763 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_762 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_761 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_760 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_759 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_758 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_757 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_756 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_755 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_754 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_753 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_752 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_751 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_750 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_749 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_748 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_747 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_746 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_745 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_744 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_743 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_742 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_741 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_740 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_739 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_738 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_737 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_736 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_735 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_734 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_733 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_732 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_731 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_730 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_729 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_728 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_727 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_726 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_725 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_724 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_723 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_722 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_721 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_720 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_719 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_718 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_717 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_716 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_715 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_714 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_713 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_712 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_711 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_710 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_709 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_708 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_707 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_706 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_705 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_704 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_703 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_702 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_701 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_700 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_699 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_698 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_697 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_696 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_695 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_694 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_693 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_692 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_691 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_690 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_689 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_688 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_687 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_686 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_685 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_684 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_683 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_682 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_681 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_680 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_679 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_678 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_677 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_676 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_675 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_674 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_673 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_672 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_671 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_669 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_668 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_666 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_665 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_663 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_662 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_657 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_656 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_655 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_654 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_653 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_651 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_650 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_649 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_648 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_647 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_645 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_644 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_643 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_642 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_641 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_640 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_639 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_638 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_637 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_635 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_626 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_625 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_624 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_623 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_621 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_620 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_618 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_617 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_616 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_615 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_614 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_612 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_611 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_609 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_608 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_606 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_605 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_604 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_603 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_602 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_600 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_599 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_598 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_597 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_596 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_595 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_594 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_593 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_592 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_591 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_590 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_589 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_588 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_587 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_586 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_585 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_584 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_583 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_582 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_581 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_580 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_579 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_578 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_577 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_576 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_575 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_574 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_573 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_572 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_570 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_569 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_567 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_566 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_565 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_563 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_561 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_560 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_559 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_558 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_557 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_556 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_555 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_554 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_551 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_549 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_548 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_547 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_546 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_545 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_543 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_542 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_537 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_536 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_534 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_533 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_531 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_530 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_529 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_527 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_524 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_522 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_521 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_520 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_518 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_517 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_512 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_510 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_509 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_507 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_506 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_505 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_504 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_503 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_501 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_500 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_499 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_498 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_497 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_496 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_495 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_494 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_493 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_492 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_491 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_490 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_489 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_488 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_487 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_486 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_485 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_484 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_483 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_482 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_481 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_480 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_479 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_478 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_477 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_476 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_474 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_473 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_472 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_471 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_470 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_467 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_465 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_464 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_463 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_462 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_461 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_459 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_458 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_457 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_455 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_453 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_452 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_451 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_450 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_449 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_448 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_447 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_446 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_445 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_443 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_441 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_440 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_438 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_437 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_435 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_434 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_431 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_429 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_428 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_426 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_425 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_424 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_423 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_422 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_419 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_416 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_413 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_411 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_410 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_409 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_408 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_407 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_405 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_404 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_402 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_401 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_400 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_399 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_398 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_397 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_396 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_395 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_394 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_393 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_392 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_391 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_390 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_389 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_388 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_387 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_386 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_385 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_384 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_383 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_382 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_381 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_380 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_379 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_378 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_377 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_376 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_375 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_374 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_371 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_369 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_368 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_367 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_366 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_365 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_364 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_363 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_362 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_359 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_357 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_356 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_354 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_353 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_351 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_350 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_349 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_348 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_347 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_345 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_344 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_341 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_340 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_339 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_338 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_337 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_336 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_335 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_333 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_332 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_331 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_330 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_329 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_327 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_326 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_320 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_317 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_315 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_314 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_313 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_308 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_307 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_306 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_305 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_303 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_302 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_301 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_300 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_299 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_297 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_296 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_295 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_294 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_293 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_292 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_291 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_290 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_289 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_288 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_287 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_286 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_285 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_284 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_283 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_282 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_281 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_280 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_279 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_278 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_277 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_276 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_275 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_273 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_272 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_271 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_270 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_269 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_267 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_266 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_265 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_263 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_261 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_260 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_258 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_257 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_256 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_255 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_254 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_251 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_249 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_248 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_246 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_245 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_244 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_243 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_242 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_240 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_237 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_236 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_235 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_234 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_233 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_232 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_231 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_230 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_219 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_212 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_210 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_209 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_208 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_207 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_206 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_203 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_201 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_200 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_199 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_198 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_197 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_195 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_194 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_193 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_192 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_191 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_190 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_189 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_188 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_187 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_186 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_184 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_183 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_182 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_181 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_180 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_179 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_177 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_176 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_175 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_174 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_172 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_171 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_169 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_167 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_165 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_164 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_162 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_161 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_159 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_155 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_153 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_152 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_150 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_149 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_148 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_147 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_146 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_145 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_141 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_138 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_136 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_135 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_134 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_133 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_131 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_129 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_128 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_126 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_125 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_123 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_122 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_121 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_119 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_116 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_114 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_113 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_111 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_110 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_109 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_104 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_102 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_101 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_100 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_99 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_98 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_97 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_96 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_95 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_94 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_93 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_92 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_91 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_90 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_89 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_88 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_87 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_86 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_85 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_84 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_83 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_82 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_81 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_80 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_79 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_78 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_77 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_76 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_75 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_74 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_73 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_71 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_70 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_68 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_67 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_66 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_65 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_64 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_63 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_62 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_61 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_59 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_58 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_56 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_55 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_53 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_52 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_51 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_50 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_49 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_47 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_46 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_43 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_42 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_41 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_40 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_39 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_38 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_37 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_35 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_34 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_32 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_31 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_30 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_29 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_28 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_27 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_26 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_25 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_23 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_22 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_20 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_19 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_17 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_16 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_15 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_14 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_13 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_11 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_10 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_8 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_7 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_5 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_4 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2221 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2218 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2215 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2185 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X4 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2173 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2170 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2143 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2140 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2137 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1936 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1930 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_1927 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1924 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1918 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1912 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1906 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_1900 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_667 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_658 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_652 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_646 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_634 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_631 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_628 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_622 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_619 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_613 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_610 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_607 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_571 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_568 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_562 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_550 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_544 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_538 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_535 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_532 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_526 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_523 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_514 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_511 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_508 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_502 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_475 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_469 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_466 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_460 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_454 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_442 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_439 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_436 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_430 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_427 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_418 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_415 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_412 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_406 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_403 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_373 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_370 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_358 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_355 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_352 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_346 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_343 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_334 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_328 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_325 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_322 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_319 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_316 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_310 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_304 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_298 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_274 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_268 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_262 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_259 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_250 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_247 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_241 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_238 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_229 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_226 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_223 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_220 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_214 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_211 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_202 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_196 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_178 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_166 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_163 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_160 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_154 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_151 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_142 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_139 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_130 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_127 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_124 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_118 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_115 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_112 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_106 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_103 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module IV_941 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_940 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_939 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_938 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_937 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_936 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_935 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_934 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_933 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_932 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_931 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_930 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_929 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_928 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_927 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_926 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_925 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_924 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_923 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_922 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_921 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_920 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_919 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_918 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_917 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_916 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_915 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_914 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_913 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_912 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_911 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_910 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_909 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_908 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_907 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_906 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_905 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_904 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_903 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_902 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_901 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_900 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_899 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_898 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_897 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_896 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_895 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_894 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_893 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_892 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_891 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_890 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_889 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_888 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_887 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_886 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_885 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_884 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_883 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_882 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_881 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_880 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_879 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_878 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_877 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_876 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_875 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_874 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_873 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_872 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_871 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_870 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_869 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_868 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_867 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_866 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_865 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_864 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_863 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_862 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_861 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_860 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_859 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_858 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_857 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_856 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_855 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_854 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_853 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_852 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_851 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_850 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_849 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_848 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_847 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_846 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_845 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_844 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_843 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_842 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_841 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_840 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_839 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_838 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_837 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_836 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_835 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_834 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_833 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_832 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_831 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_830 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_829 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_828 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_827 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_826 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_825 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_824 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_823 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_822 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_821 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_820 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_819 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_818 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_817 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_816 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_815 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_814 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_813 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_812 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_811 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_810 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_809 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_808 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_807 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_806 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_805 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_804 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_803 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_802 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_801 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_800 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_799 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_798 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_797 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_796 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_795 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_794 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_793 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_792 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_791 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_790 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_789 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_788 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_787 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_786 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_785 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_784 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_783 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_782 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_781 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_780 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_779 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_778 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_777 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_776 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_775 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_774 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_773 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_772 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_771 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_770 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_769 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_768 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_767 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_766 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_765 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_764 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_763 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_762 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_761 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_760 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_759 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_758 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_757 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_756 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_755 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_754 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_753 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_752 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_751 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_750 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_749 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_748 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_747 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_746 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_745 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_744 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_743 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_742 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_741 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_740 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_739 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_738 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_737 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_736 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_735 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_734 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_733 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_732 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_731 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_730 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_729 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_728 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_727 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_726 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_725 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_724 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_723 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_722 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_721 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_720 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_719 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_718 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_717 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_716 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_715 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_714 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_713 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_712 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_711 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_710 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_709 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_708 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_707 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_706 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_705 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_704 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_703 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_702 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_701 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_700 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_699 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_698 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_697 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_696 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_695 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_694 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_693 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_692 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_691 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_690 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_689 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_688 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_687 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_686 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_685 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_684 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_683 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_682 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_681 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_680 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_679 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_678 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_677 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_676 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_675 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_674 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_673 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_672 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_671 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_670 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_669 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_668 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_667 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_666 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_665 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_664 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_663 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_662 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_661 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_660 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_659 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_658 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_657 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_656 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_655 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_654 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_653 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_652 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_651 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_650 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_649 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_648 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_647 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_646 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_645 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_644 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_643 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_642 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_641 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_640 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_639 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_638 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_637 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_636 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_635 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_634 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_633 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_632 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_631 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_630 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_629 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_628 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_627 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_626 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_625 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_624 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_623 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_622 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_621 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_620 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_619 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_618 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_617 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_616 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_615 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_614 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_613 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_612 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_611 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_610 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_609 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_608 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_607 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_606 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_605 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_604 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_603 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_602 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_601 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_600 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_599 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_598 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_597 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_596 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_595 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_594 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_593 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_592 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_591 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_590 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_589 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_588 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_587 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_586 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_585 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_584 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_583 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_582 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_581 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_580 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_579 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_578 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_577 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_576 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_575 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_574 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_573 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_572 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_571 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_570 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_569 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_568 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_567 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_566 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_565 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_564 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_563 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_562 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_561 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_560 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_559 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_558 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_557 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_556 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_555 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_554 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_553 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_552 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_551 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_550 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_549 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_548 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_547 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_546 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_545 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_544 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_543 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_542 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_541 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_540 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_539 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_538 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_537 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_536 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_535 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_534 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_533 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_532 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_531 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_530 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_529 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_528 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_527 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_526 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_525 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_524 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_523 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_522 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_521 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_520 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_519 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_518 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_517 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_516 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_515 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_514 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_513 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_512 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_511 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_510 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_509 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_508 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_507 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_506 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_505 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_504 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_503 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_502 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_501 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_500 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_499 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_498 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_497 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_496 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_495 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_494 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_493 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_492 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_491 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_490 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_489 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_488 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_487 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_486 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_485 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_484 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_483 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_482 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_481 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_480 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_479 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_478 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_477 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_476 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_475 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_474 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_473 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_472 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_471 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_470 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_469 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_468 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_467 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_466 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_465 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_464 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_463 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_462 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_461 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_460 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_459 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_458 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_457 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_456 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_455 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_454 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_453 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_452 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_451 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_450 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_449 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_448 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_447 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_446 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_445 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_444 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_443 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_442 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_441 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_440 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_439 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_438 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_437 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_436 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_435 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_434 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_433 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_432 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_431 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_430 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_429 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_428 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_427 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_426 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_425 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_424 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_423 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_422 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_421 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_420 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_419 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_418 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_417 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_416 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_415 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_414 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_413 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_412 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_411 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_410 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_409 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_408 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_407 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_406 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_405 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_404 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_403 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_402 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_401 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_400 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_399 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_398 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_397 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_396 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_395 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_394 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_393 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_392 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_391 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_390 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_389 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_388 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_387 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_386 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_385 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_384 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_383 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_382 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_381 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_380 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_379 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_378 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_377 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_376 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_375 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_374 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_373 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_372 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_371 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_370 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_369 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_368 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_367 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_366 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_365 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_364 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_363 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_362 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_361 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_360 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_359 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_358 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_357 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_356 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_355 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_354 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_353 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_352 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_351 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_350 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_349 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_348 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_347 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_346 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_345 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_344 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_343 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_342 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_341 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_340 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_339 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_338 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_337 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_336 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_335 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_334 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_333 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_332 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_331 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_330 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_329 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_328 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_327 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_326 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_325 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_324 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_323 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_322 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_321 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_320 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_319 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_318 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_317 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_316 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_315 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_314 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_313 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_312 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_311 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_310 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_309 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_308 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_307 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_306 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_305 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_304 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_303 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_302 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_301 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_300 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_299 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_298 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_297 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_296 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_295 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_294 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_293 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_292 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_291 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_290 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_289 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_288 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_287 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_286 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_285 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_284 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_283 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_282 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_281 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_280 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_279 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_278 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_277 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_276 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_275 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_274 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_273 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_272 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_271 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_270 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_269 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_268 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_267 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_266 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_265 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_264 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_263 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_262 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_261 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_260 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_259 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_258 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_257 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_256 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_255 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_254 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_253 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_252 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_251 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_250 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_249 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_248 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_247 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_246 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_245 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_244 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_243 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_242 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_241 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_240 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_239 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_238 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_237 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_236 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_235 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_234 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_233 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_232 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_231 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_230 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_229 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_228 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_227 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_226 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_225 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_224 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_223 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_222 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_221 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_220 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_219 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_218 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_217 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_216 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_215 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_214 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_213 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_212 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_211 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_210 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_209 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_208 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_207 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_206 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_205 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_204 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_203 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_202 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_201 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_200 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_199 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_198 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_197 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_196 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_195 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_194 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_193 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_192 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_191 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_190 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_189 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_188 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_187 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_186 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_185 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_184 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_183 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_182 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_181 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_180 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_179 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_178 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_177 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_176 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_175 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_174 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_173 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_172 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_171 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_170 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_169 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_168 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_167 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_166 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_165 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_164 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_163 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_162 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_161 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_160 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_159 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_158 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_157 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_156 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_155 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_154 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_153 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_152 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_151 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_150 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_149 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_148 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_147 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_146 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_145 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_144 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_143 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_142 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_141 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_140 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_139 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_138 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_137 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_136 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_135 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_134 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_133 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_132 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_131 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_130 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_129 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_128 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_127 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_126 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_125 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_124 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_123 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_122 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_121 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_120 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_119 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_118 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_117 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_116 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_115 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_114 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_113 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_112 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_111 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_110 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_109 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_108 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_107 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_106 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_105 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_104 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_103 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_102 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_101 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_100 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_99 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_98 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_97 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_96 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_95 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_94 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_93 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_92 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_91 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_90 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_89 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_88 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_87 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_86 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_85 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_84 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_83 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_82 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_81 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_80 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_79 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_78 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_77 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_76 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_75 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_74 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_73 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_72 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_71 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_70 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_69 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_68 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_67 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_66 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_65 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_64 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_63 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_62 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_61 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_60 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_59 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_58 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_57 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_56 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_55 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_54 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_53 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_52 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_51 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_50 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_49 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_48 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_47 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_46 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_45 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_44 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_43 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_42 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_41 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_40 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_39 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_38 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_37 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_36 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_35 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_34 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_33 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_32 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_31 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_30 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_29 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_28 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_27 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_26 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_25 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_24 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_23 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_22 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_21 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_20 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_19 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_18 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_17 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_16 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_15 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_14 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_13 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_12 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_11 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_10 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_9 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_8 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_7 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_6 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_5 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_4 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_3 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_2 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module IV_1 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_N32_8 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_512 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_511 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_510 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_509 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_508 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_507 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_506 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_505 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_504 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_503 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_502 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_501 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_500 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_499 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_498 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_497 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_496 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_495 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_494 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_493 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_492 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_491 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_490 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_489 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_488 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_487 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_486 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_485 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_484 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_483 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_482 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_481 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n4) );
  BUF_X1 U2 ( .A(n3), .Z(n5) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_4 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n6, n7, n8, n9;
  assign n6 = S;

  MUX21_384 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n7), .Y(Y[0]) );
  MUX21_383 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n7), .Y(Y[1]) );
  MUX21_382 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n7), .Y(Y[2]) );
  MUX21_381 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n7), .Y(Y[3]) );
  MUX21_380 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n7), .Y(Y[4]) );
  MUX21_379 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n7), .Y(Y[5]) );
  MUX21_378 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n7), .Y(Y[6]) );
  MUX21_377 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n7), .Y(Y[7]) );
  MUX21_376 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n7), .Y(Y[8]) );
  MUX21_375 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n7), .Y(Y[9]) );
  MUX21_374 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n7), .Y(Y[10]) );
  MUX21_373 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n7), .Y(Y[11]) );
  MUX21_372 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n8), .Y(Y[12]) );
  MUX21_371 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n8), .Y(Y[13]) );
  MUX21_370 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n8), .Y(Y[14]) );
  MUX21_369 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n8), .Y(Y[15]) );
  MUX21_368 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n8), .Y(Y[16]) );
  MUX21_367 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n8), .Y(Y[17]) );
  MUX21_366 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n8), .Y(Y[18]) );
  MUX21_365 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n8), .Y(Y[19]) );
  MUX21_364 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n8), .Y(Y[20]) );
  MUX21_363 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n8), .Y(Y[21]) );
  MUX21_362 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n8), .Y(Y[22]) );
  MUX21_361 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n8), .Y(Y[23]) );
  MUX21_360 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n9), .Y(Y[24]) );
  MUX21_359 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n9), .Y(Y[25]) );
  MUX21_358 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n9), .Y(Y[26]) );
  MUX21_357 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n9), .Y(Y[27]) );
  MUX21_356 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n9), .Y(Y[28]) );
  MUX21_355 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n9), .Y(Y[29]) );
  MUX21_354 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n9), .Y(Y[30]) );
  MUX21_353 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n9), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n6), .Z(n7) );
  BUF_X1 U2 ( .A(n6), .Z(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n9) );
endmodule


module MUX21_GENERIC_N32_3 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n6, n7, n8, n9;
  assign n6 = S;

  MUX21_352 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n7), .Y(Y[0]) );
  MUX21_351 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n7), .Y(Y[1]) );
  MUX21_350 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n7), .Y(Y[2]) );
  MUX21_349 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n7), .Y(Y[3]) );
  MUX21_348 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n7), .Y(Y[4]) );
  MUX21_347 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n7), .Y(Y[5]) );
  MUX21_346 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n7), .Y(Y[6]) );
  MUX21_345 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n7), .Y(Y[7]) );
  MUX21_344 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n7), .Y(Y[8]) );
  MUX21_343 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n7), .Y(Y[9]) );
  MUX21_342 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n7), .Y(Y[10]) );
  MUX21_341 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n7), .Y(Y[11]) );
  MUX21_340 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n8), .Y(Y[12]) );
  MUX21_339 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n8), .Y(Y[13]) );
  MUX21_338 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n8), .Y(Y[14]) );
  MUX21_337 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n8), .Y(Y[15]) );
  MUX21_336 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n8), .Y(Y[16]) );
  MUX21_335 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n8), .Y(Y[17]) );
  MUX21_334 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n8), .Y(Y[18]) );
  MUX21_333 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n8), .Y(Y[19]) );
  MUX21_332 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n8), .Y(Y[20]) );
  MUX21_331 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n8), .Y(Y[21]) );
  MUX21_330 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n8), .Y(Y[22]) );
  MUX21_329 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n8), .Y(Y[23]) );
  MUX21_328 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n9), .Y(Y[24]) );
  MUX21_327 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n9), .Y(Y[25]) );
  MUX21_326 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n9), .Y(Y[26]) );
  MUX21_325 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n9), .Y(Y[27]) );
  MUX21_324 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n9), .Y(Y[28]) );
  MUX21_323 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n9), .Y(Y[29]) );
  MUX21_322 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n9), .Y(Y[30]) );
  MUX21_321 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n9), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n6), .Z(n7) );
  BUF_X1 U2 ( .A(n6), .Z(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n9) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12, n13, n14, n15, n16, n17, n18, n19;

  BUF_X1 U1 ( .A(B), .Z(n11) );
  XNOR2_X1 U2 ( .A(n12), .B(n14), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(n11), .ZN(n12) );
  CLKBUF_X1 U4 ( .A(A), .Z(n13) );
  BUF_X1 U5 ( .A(Ci), .Z(n14) );
  NAND2_X1 U6 ( .A1(n11), .A2(n13), .ZN(n19) );
  INV_X1 U7 ( .A(A), .ZN(n16) );
  INV_X1 U8 ( .A(B), .ZN(n15) );
  NAND2_X1 U9 ( .A1(n16), .A2(n15), .ZN(n17) );
  NAND2_X1 U10 ( .A1(Ci), .A2(n17), .ZN(n18) );
  NAND2_X1 U11 ( .A1(n18), .A2(n19), .ZN(Co) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  INV_X1 U1 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n7) );
  OAI21_X1 U3 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  NOR2_X1 U4 ( .A1(B), .A2(A), .ZN(n9) );
  FA_X1 U5 ( .A(A), .B(Ci), .CI(B), .S(S) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  INV_X1 U1 ( .A(n8), .ZN(n11) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n10) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n9), .ZN(S) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n9), .ZN(S) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n9), .ZN(S) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n9), .ZN(S) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n9), .ZN(S) );
endmodule


module RCA_gen_N4_101 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_404 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_403 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_402 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_401 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_100 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_400 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_399 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_398 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_397 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_99 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_396 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_395 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_394 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_393 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_98 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_392 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_391 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_390 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_389 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_97 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_388 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_387 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_386 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_385 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net181711, n7, n8, n9, n10;
  assign Co = net181711;

  XNOR2_X1 U1 ( .A(A), .B(Ci), .ZN(n10) );
  OAI21_X1 U2 ( .B1(n7), .B2(n8), .A(n9), .ZN(net181711) );
  NAND2_X1 U3 ( .A1(A), .A2(Ci), .ZN(n9) );
  NOR2_X1 U4 ( .A1(A), .A2(Ci), .ZN(n8) );
  XNOR2_X1 U5 ( .A(B), .B(n10), .ZN(S) );
  INV_X1 U6 ( .A(B), .ZN(n7) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  BUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XOR2_X1 U2 ( .A(n9), .B(n10), .Z(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U4 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XOR2_X1 U1 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(n9), .Z(n7) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n9) );
  XOR2_X1 U3 ( .A(n7), .B(n10), .Z(S) );
  OAI21_X1 U4 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U5 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(n8), .B(Ci), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(B), .Z(n7) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n9) );
  XOR2_X1 U3 ( .A(n9), .B(n10), .Z(S) );
  OAI21_X1 U4 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U5 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U6 ( .A1(A), .A2(n7), .ZN(n8) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n11), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U6 ( .A(n9), .ZN(n13) );
  XNOR2_X1 U7 ( .A(n13), .B(n12), .ZN(S) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  INV_X1 U1 ( .A(Ci), .ZN(n8) );
  NOR2_X1 U2 ( .A1(B), .A2(A), .ZN(n9) );
  OAI21_X1 U3 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  FA_X1 U5 ( .A(B), .B(A), .CI(Ci), .S(S) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(B), .Z(n7) );
  INV_X1 U2 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n8) );
  OAI21_X1 U4 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  NOR2_X1 U5 ( .A1(B), .A2(A), .ZN(n10) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n7), .S(S) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14, n15;

  CLKBUF_X1 U1 ( .A(n12), .Z(n10) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n11) );
  INV_X1 U3 ( .A(n10), .ZN(n15) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n14) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n12), .ZN(n13) );
  NAND2_X1 U7 ( .A1(n13), .A2(n14), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n11), .B(n15), .ZN(S) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(B), .Z(n9) );
  CLKBUF_X1 U2 ( .A(n14), .Z(n10) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(n9), .ZN(n13) );
  INV_X1 U5 ( .A(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n14), .ZN(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  CLKBUF_X1 U1 ( .A(n10), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n11), .Z(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n10) );
  INV_X1 U5 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n9) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n11), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U6 ( .A(n9), .ZN(n13) );
  XNOR2_X1 U7 ( .A(n13), .B(n12), .ZN(S) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n11), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U6 ( .A(n9), .ZN(n13) );
  XNOR2_X1 U7 ( .A(n13), .B(n12), .ZN(S) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(Ci), .B(n12), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(n9), .B(n13), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U5 ( .A(n13), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n12), .A2(n11), .ZN(Co) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n13) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n9) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  BUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net181054, n9, n10, n11, n12, n13;
  assign Co = net181054;

  NAND2_X1 U1 ( .A1(Ci), .A2(n12), .ZN(n11) );
  NAND2_X1 U2 ( .A1(n11), .A2(n10), .ZN(net181054) );
  INV_X1 U3 ( .A(n9), .ZN(n12) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(n13) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n9) );
  XNOR2_X1 U6 ( .A(n13), .B(n9), .ZN(S) );
  NAND2_X1 U7 ( .A1(A), .A2(B), .ZN(n10) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14, n15;

  INV_X1 U1 ( .A(A), .ZN(n10) );
  INV_X1 U2 ( .A(n9), .ZN(n15) );
  XNOR2_X1 U3 ( .A(B), .B(n10), .ZN(n9) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(n11) );
  CLKBUF_X1 U5 ( .A(B), .Z(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(A), .ZN(n14) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n9), .ZN(n13) );
  NAND2_X1 U8 ( .A1(n13), .A2(n14), .ZN(Co) );
  XNOR2_X1 U9 ( .A(n11), .B(n15), .ZN(S) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(n9), .B(n13), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U5 ( .A(n13), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n11), .A2(n12), .ZN(Co) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  INV_X1 U1 ( .A(A), .ZN(n9) );
  XNOR2_X1 U2 ( .A(B), .B(n9), .ZN(n11) );
  INV_X1 U3 ( .A(n11), .ZN(n14) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(n10) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n13) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n10), .B(n14), .ZN(S) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n10) );
  XNOR2_X1 U6 ( .A(n10), .B(n9), .ZN(S) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(B), .Z(n9) );
  INV_X1 U2 ( .A(n10), .ZN(n13) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(n9), .ZN(n12) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  INV_X1 U1 ( .A(n9), .ZN(n12) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n9) );
  XNOR2_X1 U3 ( .A(Ci), .B(n12), .ZN(S) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n11) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  AND2_X1 U1 ( .A1(A), .A2(B), .ZN(n9) );
  AOI21_X1 U2 ( .B1(Ci), .B2(n12), .A(n9), .ZN(n10) );
  INV_X1 U3 ( .A(n10), .ZN(Co) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(n11) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n13) );
  INV_X1 U6 ( .A(n13), .ZN(n12) );
  XNOR2_X1 U7 ( .A(n11), .B(n13), .ZN(S) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(n9), .B(n13), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U5 ( .A(n13), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n11), .A2(n12), .ZN(Co) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(B), .Z(n9) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(n9), .ZN(n13) );
  INV_X1 U5 ( .A(n14), .ZN(n11) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n10), .B(n14), .ZN(S) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(n10), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n10) );
  INV_X1 U4 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n9) );
  INV_X1 U6 ( .A(n8), .ZN(n12) );
  XNOR2_X1 U7 ( .A(n12), .B(n11), .ZN(S) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module RCA_gen_N4_123 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_492 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_491 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_490 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_489 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_121 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_484 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_483 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_482 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_481 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_119 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_476 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_475 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_474 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_473 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_117 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_468 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_467 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_466 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_465 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_115 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_460 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_459 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_458 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_457 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_113 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_452 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_451 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_450 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_449 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_103 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_412 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_411 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_410 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_409 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_83 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_332 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_331 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_330 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_329 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_81 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_324 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_323 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_322 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_321 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_67 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_268 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_267 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_266 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_265 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_65 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_260 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_259 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_258 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_257 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_49 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_196 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_195 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_194 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_193 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_522 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_521 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_516 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_515 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_514 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_513 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  OR2_X1 U2 ( .A1(n9), .A2(n12), .ZN(n10) );
  INV_X1 U3 ( .A(n8), .ZN(n9) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n8) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(n8), .B(Ci), .Z(S) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n10) );
  NAND2_X1 U4 ( .A1(n8), .A2(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  INV_X1 U1 ( .A(n8), .ZN(n11) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n8) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n10) );
  NAND2_X1 U4 ( .A1(n8), .A2(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(n8), .B(n12), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U5 ( .A(n12), .ZN(n9) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U7 ( .A1(n11), .A2(n10), .ZN(Co) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n8) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12, n13;

  BUF_X1 U1 ( .A(n13), .Z(n8) );
  CLKBUF_X1 U2 ( .A(B), .Z(n9) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(n9), .ZN(n12) );
  INV_X1 U5 ( .A(n13), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n8), .B(Ci), .ZN(S) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  CLKBUF_X1 U2 ( .A(n13), .Z(n9) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(n8), .ZN(n12) );
  INV_X1 U5 ( .A(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n13), .Z(n8) );
  CLKBUF_X1 U2 ( .A(B), .Z(n9) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(n9), .ZN(n12) );
  INV_X1 U5 ( .A(n8), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  BUF_X1 U1 ( .A(n12), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n11), .B(Ci), .ZN(S) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n8), .A2(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n11), .B(Ci), .ZN(S) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n8), .A2(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n11), .B(Ci), .ZN(S) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n8), .A2(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n7) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n10) );
  XNOR2_X1 U6 ( .A(n10), .B(n9), .ZN(S) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n7) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n9), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module RCA_gen_N4_124 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_496 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_495 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_494 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_493 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_122 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_488 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_487 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_486 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_485 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_120 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_480 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_479 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_478 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_477 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_118 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_472 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_471 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_470 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_469 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_116 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_464 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_463 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_462 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_461 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_114 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_456 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_455 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_454 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_453 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_104 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_416 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_415 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_414 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_413 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_84 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_336 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_335 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_334 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_333 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_82 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_328 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_327 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_326 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_325 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_68 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_272 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_271 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_270 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_269 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_66 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_264 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_263 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_262 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_261 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_200 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_199 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_198 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_197 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_40 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_160 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_159 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_158 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_157 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_34 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_136 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_135 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_134 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_133 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_128 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_124 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_123 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_122 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_121 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSAdd_N4_62 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_124 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_123 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_62 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_61 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_122 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_121 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_61 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_60 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_120 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_119 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_60 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_59 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_118 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_117 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_59 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_58 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_116 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_115 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_58 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_57 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_114 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_113 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_57 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_41 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_82 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_81 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_41 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_33 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_66 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_65 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_33 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XOR2_X1 U3 ( .A(n9), .B(n10), .Z(S) );
  INV_X1 U4 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n8) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module RCA_gen_N4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_100 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_99 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_98 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_97 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(n8), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n12), .B(Ci), .ZN(S) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(n12), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(Ci), .ZN(S) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  BUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  CLKBUF_X1 U2 ( .A(n14), .Z(n10) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n13) );
  INV_X1 U5 ( .A(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n9), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n14), .ZN(S) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  CLKBUF_X1 U2 ( .A(B), .Z(n10) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(n10), .ZN(n13) );
  INV_X1 U5 ( .A(n14), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n9), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n14), .ZN(S) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net226571, net226573, net239963, n9, n10;

  XNOR2_X1 U1 ( .A(Ci), .B(n9), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(net239963) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U4 ( .A(n9), .ZN(net226573) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net226571) );
  NAND2_X1 U6 ( .A1(net239963), .A2(net226573), .ZN(n10) );
  NAND2_X1 U7 ( .A1(net226571), .A2(n10), .ZN(Co) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  OR2_X1 U2 ( .A1(n10), .A2(n13), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  OR2_X1 U2 ( .A1(n10), .A2(n13), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  OR2_X1 U2 ( .A1(n10), .A2(n13), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  OR2_X1 U2 ( .A1(n10), .A2(n13), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net225330, net225331, net239344, net240011, n9;

  XNOR2_X1 U1 ( .A(Ci), .B(n9), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(net240011) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n9) );
  OR2_X1 U4 ( .A1(net239344), .A2(n9), .ZN(net225331) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net225330) );
  INV_X1 U6 ( .A(net240011), .ZN(net239344) );
  NAND2_X1 U7 ( .A1(net225330), .A2(net225331), .ZN(Co) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(n14), .Z(n9) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n13) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n14), .ZN(S) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(n14), .Z(n9) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n13) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n14), .B(Ci), .ZN(S) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net223696, net223698, net241961, net242957, n9, n10;

  XNOR2_X1 U1 ( .A(Ci), .B(n9), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(net241961) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n9) );
  CLKBUF_X1 U4 ( .A(n9), .Z(net242957) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net223696) );
  INV_X1 U6 ( .A(net242957), .ZN(net223698) );
  NAND2_X1 U7 ( .A1(net241961), .A2(net223698), .ZN(n10) );
  NAND2_X1 U8 ( .A1(net223696), .A2(n10), .ZN(Co) );
endmodule


module MUX21_941 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_941 UIV ( .A(S), .Y(SB) );
  ND2_2823 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2822 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2821 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_940 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_940 UIV ( .A(S), .Y(SB) );
  ND2_2820 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2819 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2818 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_939 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_939 UIV ( .A(S), .Y(SB) );
  ND2_2817 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2816 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2815 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_938 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_938 UIV ( .A(S), .Y(SB) );
  ND2_2814 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2813 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2812 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_937 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_937 UIV ( .A(S), .Y(SB) );
  ND2_2811 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2810 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2809 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_936 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_936 UIV ( .A(S), .Y(SB) );
  ND2_2808 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2807 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2806 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_935 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_935 UIV ( .A(S), .Y(SB) );
  ND2_2805 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2804 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2803 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_934 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_934 UIV ( .A(S), .Y(SB) );
  ND2_2802 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2801 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2800 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_933 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_933 UIV ( .A(S), .Y(SB) );
  ND2_2799 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2798 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2797 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_932 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_932 UIV ( .A(S), .Y(SB) );
  ND2_2796 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2795 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2794 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_908 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_908 UIV ( .A(S), .Y(SB) );
  ND2_2724 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2723 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2722 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_907 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_907 UIV ( .A(S), .Y(SB) );
  ND2_2721 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2720 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2719 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_906 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_906 UIV ( .A(S), .Y(SB) );
  ND2_2718 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2717 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2716 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_905 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_905 UIV ( .A(S), .Y(SB) );
  ND2_2715 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2714 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2713 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_904 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_904 UIV ( .A(S), .Y(SB) );
  ND2_2712 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2711 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2710 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_912 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_912 UIV ( .A(S), .Y(SB) );
  ND2_2736 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2735 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2734 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_911 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_911 UIV ( .A(S), .Y(SB) );
  ND2_2733 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2732 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2731 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_910 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_910 UIV ( .A(S), .Y(SB) );
  ND2_2730 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2729 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2728 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_909 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_909 UIV ( .A(S), .Y(SB) );
  ND2_2727 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2726 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2725 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_576 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_576 UIV ( .A(S), .Y(SB) );
  ND2_1728 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1727 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1726 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_575 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_575 UIV ( .A(S), .Y(SB) );
  ND2_1725 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1724 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1723 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_574 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_574 UIV ( .A(S), .Y(SB) );
  ND2_1722 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1721 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1720 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_573 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_573 UIV ( .A(S), .Y(SB) );
  ND2_1719 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1718 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1717 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_572 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_572 UIV ( .A(S), .Y(SB) );
  ND2_1716 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1715 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1714 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_571 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_571 UIV ( .A(S), .Y(SB) );
  ND2_1713 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1712 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1711 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_570 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_570 UIV ( .A(S), .Y(SB) );
  ND2_1710 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1709 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1708 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_569 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_569 UIV ( .A(S), .Y(SB) );
  ND2_1707 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1706 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1705 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_568 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_568 UIV ( .A(S), .Y(SB) );
  ND2_1704 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1703 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1702 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_567 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_567 UIV ( .A(S), .Y(SB) );
  ND2_1701 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1700 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1699 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_566 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_566 UIV ( .A(S), .Y(SB) );
  ND2_1698 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1697 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1696 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_565 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_565 UIV ( .A(S), .Y(SB) );
  ND2_1695 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1694 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1693 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_564 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_564 UIV ( .A(S), .Y(SB) );
  ND2_1692 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1691 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1690 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_563 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_563 UIV ( .A(S), .Y(SB) );
  ND2_1689 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1688 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1687 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_562 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_562 UIV ( .A(S), .Y(SB) );
  ND2_1686 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1685 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1684 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_561 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_561 UIV ( .A(S), .Y(SB) );
  ND2_1683 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1682 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1681 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_560 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_560 UIV ( .A(S), .Y(SB) );
  ND2_1680 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1679 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1678 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_559 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_559 UIV ( .A(S), .Y(SB) );
  ND2_1677 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1676 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1675 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_558 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_558 UIV ( .A(S), .Y(SB) );
  ND2_1674 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1673 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1672 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_557 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_557 UIV ( .A(S), .Y(SB) );
  ND2_1671 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1670 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1669 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_556 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_556 UIV ( .A(S), .Y(SB) );
  ND2_1668 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1667 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1666 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_555 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_555 UIV ( .A(S), .Y(SB) );
  ND2_1665 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1664 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1663 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_554 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_554 UIV ( .A(S), .Y(SB) );
  ND2_1662 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1661 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1660 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_553 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_553 UIV ( .A(S), .Y(SB) );
  ND2_1659 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1658 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1657 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_552 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_552 UIV ( .A(S), .Y(SB) );
  ND2_1656 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1655 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1654 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_551 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_551 UIV ( .A(S), .Y(SB) );
  ND2_1653 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1652 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1651 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_550 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_550 UIV ( .A(S), .Y(SB) );
  ND2_1650 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1649 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1648 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_549 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_549 UIV ( .A(S), .Y(SB) );
  ND2_1647 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1646 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1645 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_548 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_548 UIV ( .A(S), .Y(SB) );
  ND2_1644 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1643 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1642 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_547 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_547 UIV ( .A(S), .Y(SB) );
  ND2_1641 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1640 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1639 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_546 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_546 UIV ( .A(S), .Y(SB) );
  ND2_1638 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1637 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1636 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_545 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_545 UIV ( .A(S), .Y(SB) );
  ND2_1635 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1634 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1633 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_544 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_544 UIV ( .A(S), .Y(SB) );
  ND2_1632 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1631 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1630 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_543 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_543 UIV ( .A(S), .Y(SB) );
  ND2_1629 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1628 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1627 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_542 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_542 UIV ( .A(S), .Y(SB) );
  ND2_1626 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1625 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1624 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_541 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_541 UIV ( .A(S), .Y(SB) );
  ND2_1623 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1622 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1621 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_540 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_540 UIV ( .A(S), .Y(SB) );
  ND2_1620 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1619 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1618 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_539 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_539 UIV ( .A(S), .Y(SB) );
  ND2_1617 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1616 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1615 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_538 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_538 UIV ( .A(S), .Y(SB) );
  ND2_1614 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1613 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1612 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_537 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_537 UIV ( .A(S), .Y(SB) );
  ND2_1611 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1610 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1609 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_536 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_536 UIV ( .A(S), .Y(SB) );
  ND2_1608 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1607 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1606 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_535 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_535 UIV ( .A(S), .Y(SB) );
  ND2_1605 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1604 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1603 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_534 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_534 UIV ( .A(S), .Y(SB) );
  ND2_1602 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1601 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1600 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_533 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_533 UIV ( .A(S), .Y(SB) );
  ND2_1599 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1598 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1597 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_532 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_532 UIV ( .A(S), .Y(SB) );
  ND2_1596 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1595 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1594 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_531 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_531 UIV ( .A(S), .Y(SB) );
  ND2_1593 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1592 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1591 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_530 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_530 UIV ( .A(S), .Y(SB) );
  ND2_1590 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1589 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1588 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_529 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_529 UIV ( .A(S), .Y(SB) );
  ND2_1587 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1586 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1585 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_528 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_528 UIV ( .A(S), .Y(SB) );
  ND2_1584 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1583 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1582 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_527 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_527 UIV ( .A(S), .Y(SB) );
  ND2_1581 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1580 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1579 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_526 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_526 UIV ( .A(S), .Y(SB) );
  ND2_1578 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1577 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1576 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_525 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_525 UIV ( .A(S), .Y(SB) );
  ND2_1575 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1574 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1573 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_524 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_524 UIV ( .A(S), .Y(SB) );
  ND2_1572 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1571 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1570 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_523 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_523 UIV ( .A(S), .Y(SB) );
  ND2_1569 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1568 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1567 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_522 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_522 UIV ( .A(S), .Y(SB) );
  ND2_1566 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1565 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1564 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_521 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_521 UIV ( .A(S), .Y(SB) );
  ND2_1563 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1562 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1561 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_520 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_520 UIV ( .A(S), .Y(SB) );
  ND2_1560 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1559 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1558 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_519 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_519 UIV ( .A(S), .Y(SB) );
  ND2_1557 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1556 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1555 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_518 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_518 UIV ( .A(S), .Y(SB) );
  ND2_1554 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1553 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1552 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_517 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_517 UIV ( .A(S), .Y(SB) );
  ND2_1551 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1550 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1549 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_516 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_516 UIV ( .A(S), .Y(SB) );
  ND2_1548 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1547 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1546 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_515 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_515 UIV ( .A(S), .Y(SB) );
  ND2_1545 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1544 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1543 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_514 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_514 UIV ( .A(S), .Y(SB) );
  ND2_1542 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1541 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1540 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_513 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_513 UIV ( .A(S), .Y(SB) );
  ND2_1539 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1538 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1537 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_512 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_512 UIV ( .A(S), .Y(SB) );
  ND2_1536 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1535 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1534 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_511 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_511 UIV ( .A(S), .Y(SB) );
  ND2_1533 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1532 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1531 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_510 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_510 UIV ( .A(S), .Y(SB) );
  ND2_1530 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1529 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1528 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_509 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_509 UIV ( .A(S), .Y(SB) );
  ND2_1527 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1526 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1525 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_508 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_508 UIV ( .A(S), .Y(SB) );
  ND2_1524 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1523 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1522 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_507 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_507 UIV ( .A(S), .Y(SB) );
  ND2_1521 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1520 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1519 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_506 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_506 UIV ( .A(S), .Y(SB) );
  ND2_1518 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1517 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1516 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_505 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_505 UIV ( .A(S), .Y(SB) );
  ND2_1515 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1514 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1513 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_504 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_504 UIV ( .A(S), .Y(SB) );
  ND2_1512 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1511 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1510 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_503 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_503 UIV ( .A(S), .Y(SB) );
  ND2_1509 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1508 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1507 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_502 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_502 UIV ( .A(S), .Y(SB) );
  ND2_1506 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1505 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1504 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_501 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_501 UIV ( .A(S), .Y(SB) );
  ND2_1503 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1502 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1501 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_500 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_500 UIV ( .A(S), .Y(SB) );
  ND2_1500 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1499 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1498 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_499 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_499 UIV ( .A(S), .Y(SB) );
  ND2_1497 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1496 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1495 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_498 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_498 UIV ( .A(S), .Y(SB) );
  ND2_1494 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1493 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1492 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_497 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_497 UIV ( .A(S), .Y(SB) );
  ND2_1491 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1490 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1489 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_496 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_496 UIV ( .A(S), .Y(SB) );
  ND2_1488 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1487 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1486 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_495 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_495 UIV ( .A(S), .Y(SB) );
  ND2_1485 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1484 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1483 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_494 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_494 UIV ( .A(S), .Y(SB) );
  ND2_1482 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1481 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1480 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_493 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_493 UIV ( .A(S), .Y(SB) );
  ND2_1479 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1478 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1477 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_492 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_492 UIV ( .A(S), .Y(SB) );
  ND2_1476 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1475 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1474 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_491 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_491 UIV ( .A(S), .Y(SB) );
  ND2_1473 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1472 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1471 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_490 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_490 UIV ( .A(S), .Y(SB) );
  ND2_1470 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1469 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1468 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_489 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_489 UIV ( .A(S), .Y(SB) );
  ND2_1467 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1466 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1465 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_488 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_488 UIV ( .A(S), .Y(SB) );
  ND2_1464 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1463 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1462 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_487 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_487 UIV ( .A(S), .Y(SB) );
  ND2_1461 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1460 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1459 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_486 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_486 UIV ( .A(S), .Y(SB) );
  ND2_1458 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1457 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1456 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_485 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_485 UIV ( .A(S), .Y(SB) );
  ND2_1455 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1454 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1453 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_484 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_484 UIV ( .A(S), .Y(SB) );
  ND2_1452 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1451 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1450 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_483 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_483 UIV ( .A(S), .Y(SB) );
  ND2_1449 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1448 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1447 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_482 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_482 UIV ( .A(S), .Y(SB) );
  ND2_1446 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1445 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1444 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_481 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_481 UIV ( .A(S), .Y(SB) );
  ND2_1443 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1442 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1441 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_930 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_930 UIV ( .A(S), .Y(SB) );
  ND2_2790 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2789 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2788 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_929 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_929 UIV ( .A(S), .Y(SB) );
  ND2_2787 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2786 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2785 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_928 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_928 UIV ( .A(S), .Y(SB) );
  ND2_2784 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2783 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2782 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_927 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_927 UIV ( .A(S), .Y(SB) );
  ND2_2781 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2780 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2779 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_926 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_926 UIV ( .A(S), .Y(SB) );
  ND2_2778 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2777 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2776 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_925 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_925 UIV ( .A(S), .Y(SB) );
  ND2_2775 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2774 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2773 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_924 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_924 UIV ( .A(S), .Y(SB) );
  ND2_2772 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2771 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2770 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_923 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_923 UIV ( .A(S), .Y(SB) );
  ND2_2769 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2768 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2767 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_922 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_922 UIV ( .A(S), .Y(SB) );
  ND2_2766 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2765 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2764 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_919 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_919 UIV ( .A(S), .Y(SB) );
  ND2_2757 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2756 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2755 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_918 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_918 UIV ( .A(S), .Y(SB) );
  ND2_2754 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2753 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2752 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_917 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_917 UIV ( .A(S), .Y(SB) );
  ND2_2751 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2750 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2749 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_916 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_916 UIV ( .A(S), .Y(SB) );
  ND2_2748 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2747 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2746 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_915 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_915 UIV ( .A(S), .Y(SB) );
  ND2_2745 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2744 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2743 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_914 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_914 UIV ( .A(S), .Y(SB) );
  ND2_2742 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2741 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2740 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_903 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_903 UIV ( .A(S), .Y(SB) );
  ND2_2709 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2708 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2707 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_902 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_902 UIV ( .A(S), .Y(SB) );
  ND2_2706 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2705 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2704 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_901 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_901 UIV ( .A(S), .Y(SB) );
  ND2_2703 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2702 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2701 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_900 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_900 UIV ( .A(S), .Y(SB) );
  ND2_2700 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2699 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2698 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_899 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_899 UIV ( .A(S), .Y(SB) );
  ND2_2697 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2696 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2695 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_898 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_898 UIV ( .A(S), .Y(SB) );
  ND2_2694 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2693 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2692 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_897 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_897 UIV ( .A(S), .Y(SB) );
  ND2_2691 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2690 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2689 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_896 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_896 UIV ( .A(S), .Y(SB) );
  ND2_2688 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2687 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2686 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_895 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_895 UIV ( .A(S), .Y(SB) );
  ND2_2685 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2684 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2683 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_894 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_894 UIV ( .A(S), .Y(SB) );
  ND2_2682 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2681 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2680 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_893 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_893 UIV ( .A(S), .Y(SB) );
  ND2_2679 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2678 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2677 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_892 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_892 UIV ( .A(S), .Y(SB) );
  ND2_2676 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2675 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2674 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_891 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_891 UIV ( .A(S), .Y(SB) );
  ND2_2673 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2672 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2671 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_890 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_890 UIV ( .A(S), .Y(SB) );
  ND2_2670 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2669 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2668 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_889 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_889 UIV ( .A(S), .Y(SB) );
  ND2_2667 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2666 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2665 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_888 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_888 UIV ( .A(S), .Y(SB) );
  ND2_2664 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2663 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2662 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_855 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_855 UIV ( .A(S), .Y(SB) );
  ND2_2565 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2564 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2563 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_854 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_854 UIV ( .A(S), .Y(SB) );
  ND2_2562 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2561 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2560 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_853 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_853 UIV ( .A(S), .Y(SB) );
  ND2_2559 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2558 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2557 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_852 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_852 UIV ( .A(S), .Y(SB) );
  ND2_2556 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2555 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2554 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_851 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_851 UIV ( .A(S), .Y(SB) );
  ND2_2553 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2552 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2551 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_850 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_850 UIV ( .A(S), .Y(SB) );
  ND2_2550 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2549 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2548 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_849 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_849 UIV ( .A(S), .Y(SB) );
  ND2_2547 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2546 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2545 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_848 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_848 UIV ( .A(S), .Y(SB) );
  ND2_2544 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2543 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2542 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_847 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_847 UIV ( .A(S), .Y(SB) );
  ND2_2541 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2540 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2539 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_846 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_846 UIV ( .A(S), .Y(SB) );
  ND2_2538 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2537 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2536 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_845 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_845 UIV ( .A(S), .Y(SB) );
  ND2_2535 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2534 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2533 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_844 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_844 UIV ( .A(S), .Y(SB) );
  ND2_2532 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2531 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2530 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_843 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_843 UIV ( .A(S), .Y(SB) );
  ND2_2529 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2528 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2527 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_842 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_842 UIV ( .A(S), .Y(SB) );
  ND2_2526 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2525 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2524 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_841 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_841 UIV ( .A(S), .Y(SB) );
  ND2_2523 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2522 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2521 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_840 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_840 UIV ( .A(S), .Y(SB) );
  ND2_2520 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2519 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2518 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_839 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_839 UIV ( .A(S), .Y(SB) );
  ND2_2517 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2516 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2515 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_838 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_838 UIV ( .A(S), .Y(SB) );
  ND2_2514 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2513 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2512 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_837 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_837 UIV ( .A(S), .Y(SB) );
  ND2_2511 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2510 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2509 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_836 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_836 UIV ( .A(S), .Y(SB) );
  ND2_2508 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2507 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2506 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_835 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_835 UIV ( .A(S), .Y(SB) );
  ND2_2505 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2504 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2503 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_834 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_834 UIV ( .A(S), .Y(SB) );
  ND2_2502 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2501 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2500 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_833 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_833 UIV ( .A(S), .Y(SB) );
  ND2_2499 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2498 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2497 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_832 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_832 UIV ( .A(S), .Y(SB) );
  ND2_2496 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2495 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2494 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_831 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_831 UIV ( .A(S), .Y(SB) );
  ND2_2493 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2492 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2491 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_830 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_830 UIV ( .A(S), .Y(SB) );
  ND2_2490 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2489 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2488 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_829 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_829 UIV ( .A(S), .Y(SB) );
  ND2_2487 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2486 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2485 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_828 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_828 UIV ( .A(S), .Y(SB) );
  ND2_2484 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2483 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2482 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_827 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_827 UIV ( .A(S), .Y(SB) );
  ND2_2481 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2480 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2479 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_826 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_826 UIV ( .A(S), .Y(SB) );
  ND2_2478 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2477 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2476 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_825 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_825 UIV ( .A(S), .Y(SB) );
  ND2_2475 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2474 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2473 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_824 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_824 UIV ( .A(S), .Y(SB) );
  ND2_2472 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2471 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2470 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_823 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_823 UIV ( .A(S), .Y(SB) );
  ND2_2469 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2468 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2467 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_822 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_822 UIV ( .A(S), .Y(SB) );
  ND2_2466 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2465 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2464 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_821 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_821 UIV ( .A(S), .Y(SB) );
  ND2_2463 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2462 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2461 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_820 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_820 UIV ( .A(S), .Y(SB) );
  ND2_2460 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2459 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2458 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_819 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_819 UIV ( .A(S), .Y(SB) );
  ND2_2457 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2456 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2455 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_818 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_818 UIV ( .A(S), .Y(SB) );
  ND2_2454 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2453 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2452 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_817 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_817 UIV ( .A(S), .Y(SB) );
  ND2_2451 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2450 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2449 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_816 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_816 UIV ( .A(S), .Y(SB) );
  ND2_2448 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2447 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2446 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_815 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_815 UIV ( .A(S), .Y(SB) );
  ND2_2445 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2444 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2443 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_814 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_814 UIV ( .A(S), .Y(SB) );
  ND2_2442 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2441 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2440 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_813 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_813 UIV ( .A(S), .Y(SB) );
  ND2_2439 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2438 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2437 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_812 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_812 UIV ( .A(S), .Y(SB) );
  ND2_2436 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2435 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2434 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_811 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_811 UIV ( .A(S), .Y(SB) );
  ND2_2433 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2432 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2431 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_810 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_810 UIV ( .A(S), .Y(SB) );
  ND2_2430 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2429 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2428 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_809 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_809 UIV ( .A(S), .Y(SB) );
  ND2_2427 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2426 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2425 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_808 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_808 UIV ( .A(S), .Y(SB) );
  ND2_2424 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2423 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2422 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_807 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_807 UIV ( .A(S), .Y(SB) );
  ND2_2421 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2420 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2419 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_805 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_805 UIV ( .A(S), .Y(SB) );
  ND2_2415 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2414 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2413 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_804 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_804 UIV ( .A(S), .Y(SB) );
  ND2_2412 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2411 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2410 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_803 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_803 UIV ( .A(S), .Y(SB) );
  ND2_2409 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2408 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2407 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_802 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_802 UIV ( .A(S), .Y(SB) );
  ND2_2406 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2405 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2404 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_801 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_801 UIV ( .A(S), .Y(SB) );
  ND2_2403 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2402 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2401 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_800 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_800 UIV ( .A(S), .Y(SB) );
  ND2_2400 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2399 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2398 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_799 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_799 UIV ( .A(S), .Y(SB) );
  ND2_2397 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2396 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2395 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_797 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_797 UIV ( .A(S), .Y(SB) );
  ND2_2391 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2390 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2389 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_796 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_796 UIV ( .A(S), .Y(SB) );
  ND2_2388 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2387 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2386 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_795 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_795 UIV ( .A(S), .Y(SB) );
  ND2_2385 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2384 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2383 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_794 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_794 UIV ( .A(S), .Y(SB) );
  ND2_2382 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2381 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2380 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_793 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_793 UIV ( .A(S), .Y(SB) );
  ND2_2379 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2378 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2377 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_792 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_792 UIV ( .A(S), .Y(SB) );
  ND2_2376 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2375 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2374 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_791 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_791 UIV ( .A(S), .Y(SB) );
  ND2_2373 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2372 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2371 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_790 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_790 UIV ( .A(S), .Y(SB) );
  ND2_2370 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2369 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2368 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_789 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_789 UIV ( .A(S), .Y(SB) );
  ND2_2367 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2366 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2365 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_788 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_788 UIV ( .A(S), .Y(SB) );
  ND2_2364 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2363 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2362 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_787 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_787 UIV ( .A(S), .Y(SB) );
  ND2_2361 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2360 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2359 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_786 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_786 UIV ( .A(S), .Y(SB) );
  ND2_2358 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2357 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2356 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_785 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_785 UIV ( .A(S), .Y(SB) );
  ND2_2355 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2354 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2353 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_784 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_784 UIV ( .A(S), .Y(SB) );
  ND2_2352 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2351 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2350 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_783 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_783 UIV ( .A(S), .Y(SB) );
  ND2_2349 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2348 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2347 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_782 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_782 UIV ( .A(S), .Y(SB) );
  ND2_2346 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2345 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2344 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_781 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_781 UIV ( .A(S), .Y(SB) );
  ND2_2343 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2342 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2341 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_780 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_780 UIV ( .A(S), .Y(SB) );
  ND2_2340 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2339 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2338 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_779 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_779 UIV ( .A(S), .Y(SB) );
  ND2_2337 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2336 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2335 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_778 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_778 UIV ( .A(S), .Y(SB) );
  ND2_2334 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2333 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2332 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_777 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_777 UIV ( .A(S), .Y(SB) );
  ND2_2331 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2330 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2329 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_776 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_776 UIV ( .A(S), .Y(SB) );
  ND2_2328 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2327 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2326 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_775 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_775 UIV ( .A(S), .Y(SB) );
  ND2_2325 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2324 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2323 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_774 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_774 UIV ( .A(S), .Y(SB) );
  ND2_2322 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2321 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2320 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_773 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_773 UIV ( .A(S), .Y(SB) );
  ND2_2319 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2318 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2317 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_772 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_772 UIV ( .A(S), .Y(SB) );
  ND2_2316 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2315 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2314 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_771 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_771 UIV ( .A(S), .Y(SB) );
  ND2_2313 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2312 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2311 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_768 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_768 UIV ( .A(S), .Y(SB) );
  ND2_2304 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2303 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2302 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_767 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_767 UIV ( .A(S), .Y(SB) );
  ND2_2301 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2300 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2299 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_766 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_766 UIV ( .A(S), .Y(SB) );
  ND2_2298 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2297 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2296 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_765 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_765 UIV ( .A(S), .Y(SB) );
  ND2_2295 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2294 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2293 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_764 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_764 UIV ( .A(S), .Y(SB) );
  ND2_2292 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2291 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2290 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_763 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_763 UIV ( .A(S), .Y(SB) );
  ND2_2289 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2288 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2287 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_762 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_762 UIV ( .A(S), .Y(SB) );
  ND2_2286 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2285 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2284 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_761 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_761 UIV ( .A(S), .Y(SB) );
  ND2_2283 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2282 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2281 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_760 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_760 UIV ( .A(S), .Y(SB) );
  ND2_2280 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2279 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2278 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_759 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_759 UIV ( .A(S), .Y(SB) );
  ND2_2277 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2276 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2275 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_758 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_758 UIV ( .A(S), .Y(SB) );
  ND2_2274 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2273 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2272 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_757 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_757 UIV ( .A(S), .Y(SB) );
  ND2_2271 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2270 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2269 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_756 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_756 UIV ( .A(S), .Y(SB) );
  ND2_2268 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2267 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2266 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_755 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_755 UIV ( .A(S), .Y(SB) );
  ND2_2265 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2264 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2263 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_754 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_754 UIV ( .A(S), .Y(SB) );
  ND2_2262 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2261 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2260 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_753 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_753 UIV ( .A(S), .Y(SB) );
  ND2_2259 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2258 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2257 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_752 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_752 UIV ( .A(S), .Y(SB) );
  ND2_2256 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2255 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2254 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_751 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_751 UIV ( .A(S), .Y(SB) );
  ND2_2253 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2252 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2251 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_750 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_750 UIV ( .A(S), .Y(SB) );
  ND2_2250 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2249 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2248 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_749 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_749 UIV ( .A(S), .Y(SB) );
  ND2_2247 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2246 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2245 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_748 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_748 UIV ( .A(S), .Y(SB) );
  ND2_2244 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2243 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2242 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_747 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_747 UIV ( .A(S), .Y(SB) );
  ND2_2241 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2240 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2239 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_746 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_746 UIV ( .A(S), .Y(SB) );
  ND2_2238 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2237 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2236 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_745 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_745 UIV ( .A(S), .Y(SB) );
  ND2_2235 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2234 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2233 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_744 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_744 UIV ( .A(S), .Y(SB) );
  ND2_2232 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2231 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2230 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_738 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_738 UIV ( .A(S), .Y(SB) );
  ND2_2214 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2213 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2212 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_737 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_737 UIV ( .A(S), .Y(SB) );
  ND2_2211 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2210 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2209 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_736 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_736 UIV ( .A(S), .Y(SB) );
  ND2_2208 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2207 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2206 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_734 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_734 UIV ( .A(S), .Y(SB) );
  ND2_2202 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2201 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2200 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_733 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_733 UIV ( .A(S), .Y(SB) );
  ND2_2199 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2198 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2197 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_731 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_731 UIV ( .A(S), .Y(SB) );
  ND2_2193 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2192 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2191 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_730 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_730 UIV ( .A(S), .Y(SB) );
  ND2_2190 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2189 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2188 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_728 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_728 UIV ( .A(S), .Y(SB) );
  ND2_2184 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2183 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2182 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_727 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_727 UIV ( .A(S), .Y(SB) );
  ND2_2181 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2180 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2179 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_726 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_726 UIV ( .A(S), .Y(SB) );
  ND2_2178 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2177 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2176 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_723 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_723 UIV ( .A(S), .Y(SB) );
  ND2_2169 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2168 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2167 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_722 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_722 UIV ( .A(S), .Y(SB) );
  ND2_2166 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2165 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2164 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_721 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_721 UIV ( .A(S), .Y(SB) );
  ND2_2163 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2162 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2161 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_720 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_720 UIV ( .A(S), .Y(SB) );
  ND2_2160 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2159 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2158 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_719 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_719 UIV ( .A(S), .Y(SB) );
  ND2_2157 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2156 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2155 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_718 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_718 UIV ( .A(S), .Y(SB) );
  ND2_2154 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2153 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2152 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_717 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_717 UIV ( .A(S), .Y(SB) );
  ND2_2151 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2150 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2149 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_716 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_716 UIV ( .A(S), .Y(SB) );
  ND2_2148 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2147 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2146 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_712 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_712 UIV ( .A(S), .Y(SB) );
  ND2_2136 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2135 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2134 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_710 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_710 UIV ( .A(S), .Y(SB) );
  ND2_2130 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2129 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2128 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_708 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_708 UIV ( .A(S), .Y(SB) );
  ND2_2124 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2123 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2122 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_707 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_707 UIV ( .A(S), .Y(SB) );
  ND2_2121 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2120 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2119 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_706 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_706 UIV ( .A(S), .Y(SB) );
  ND2_2118 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2117 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2116 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_705 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_705 UIV ( .A(S), .Y(SB) );
  ND2_2115 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2114 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2113 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_704 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_704 UIV ( .A(S), .Y(SB) );
  ND2_2112 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2111 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2110 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_703 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_703 UIV ( .A(S), .Y(SB) );
  ND2_2109 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2108 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2107 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_702 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_702 UIV ( .A(S), .Y(SB) );
  ND2_2106 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2105 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2104 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_701 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_701 UIV ( .A(S), .Y(SB) );
  ND2_2103 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2102 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2101 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_700 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_700 UIV ( .A(S), .Y(SB) );
  ND2_2100 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2099 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2098 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_699 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_699 UIV ( .A(S), .Y(SB) );
  ND2_2097 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2096 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2095 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_698 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_698 UIV ( .A(S), .Y(SB) );
  ND2_2094 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2093 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2092 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_697 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_697 UIV ( .A(S), .Y(SB) );
  ND2_2091 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2090 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2089 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_696 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_696 UIV ( .A(S), .Y(SB) );
  ND2_2088 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2087 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2086 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_695 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_695 UIV ( .A(S), .Y(SB) );
  ND2_2085 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2084 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2083 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_694 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_694 UIV ( .A(S), .Y(SB) );
  ND2_2082 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2081 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2080 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_693 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_693 UIV ( .A(S), .Y(SB) );
  ND2_2079 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2078 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2077 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_692 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_692 UIV ( .A(S), .Y(SB) );
  ND2_2076 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2075 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2074 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_691 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_691 UIV ( .A(S), .Y(SB) );
  ND2_2073 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2072 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2071 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_690 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_690 UIV ( .A(S), .Y(SB) );
  ND2_2070 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2069 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2068 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_689 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_689 UIV ( .A(S), .Y(SB) );
  ND2_2067 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2066 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2065 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_688 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_688 UIV ( .A(S), .Y(SB) );
  ND2_2064 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2063 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2062 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_687 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_687 UIV ( .A(S), .Y(SB) );
  ND2_2061 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2060 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2059 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_686 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_686 UIV ( .A(S), .Y(SB) );
  ND2_2058 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2057 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2056 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_685 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_685 UIV ( .A(S), .Y(SB) );
  ND2_2055 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2054 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2053 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_684 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_684 UIV ( .A(S), .Y(SB) );
  ND2_2052 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2051 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2050 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_683 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_683 UIV ( .A(S), .Y(SB) );
  ND2_2049 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2048 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2047 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_682 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_682 UIV ( .A(S), .Y(SB) );
  ND2_2046 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2045 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2044 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_681 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_681 UIV ( .A(S), .Y(SB) );
  ND2_2043 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2042 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2041 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_680 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_680 UIV ( .A(S), .Y(SB) );
  ND2_2040 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2039 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2038 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_679 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_679 UIV ( .A(S), .Y(SB) );
  ND2_2037 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2036 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2035 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_678 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_678 UIV ( .A(S), .Y(SB) );
  ND2_2034 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2033 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2032 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_677 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_677 UIV ( .A(S), .Y(SB) );
  ND2_2031 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2030 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2029 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_676 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_676 UIV ( .A(S), .Y(SB) );
  ND2_2028 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2027 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2026 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_675 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_675 UIV ( .A(S), .Y(SB) );
  ND2_2025 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2024 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2023 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_674 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_674 UIV ( .A(S), .Y(SB) );
  ND2_2022 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2021 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2020 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_673 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_673 UIV ( .A(S), .Y(SB) );
  ND2_2019 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2018 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2017 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_672 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_672 UIV ( .A(S), .Y(SB) );
  ND2_2016 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2015 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2014 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_671 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_671 UIV ( .A(S), .Y(SB) );
  ND2_2013 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2012 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2011 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_670 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_670 UIV ( .A(S), .Y(SB) );
  ND2_2010 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2009 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2008 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_669 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_669 UIV ( .A(S), .Y(SB) );
  ND2_2007 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2006 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2005 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_668 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_668 UIV ( .A(S), .Y(SB) );
  ND2_2004 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2003 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2002 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_667 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_667 UIV ( .A(S), .Y(SB) );
  ND2_2001 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2000 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1999 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_666 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_666 UIV ( .A(S), .Y(SB) );
  ND2_1998 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1997 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1996 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_665 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_665 UIV ( .A(S), .Y(SB) );
  ND2_1995 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1994 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1993 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_664 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_664 UIV ( .A(S), .Y(SB) );
  ND2_1992 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1991 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1990 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_663 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_663 UIV ( .A(S), .Y(SB) );
  ND2_1989 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1988 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1987 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_662 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_662 UIV ( .A(S), .Y(SB) );
  ND2_1986 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1985 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1984 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_661 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_661 UIV ( .A(S), .Y(SB) );
  ND2_1983 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1982 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1981 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_660 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_660 UIV ( .A(S), .Y(SB) );
  ND2_1980 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1979 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1978 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_659 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_659 UIV ( .A(S), .Y(SB) );
  ND2_1977 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1976 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1975 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_658 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_658 UIV ( .A(S), .Y(SB) );
  ND2_1974 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1973 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1972 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_657 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_657 UIV ( .A(S), .Y(SB) );
  ND2_1971 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1970 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1969 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_656 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_656 UIV ( .A(S), .Y(SB) );
  ND2_1968 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1967 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1966 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_655 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_655 UIV ( .A(S), .Y(SB) );
  ND2_1965 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1964 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1963 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_654 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_654 UIV ( .A(S), .Y(SB) );
  ND2_1962 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1961 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1960 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_653 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_653 UIV ( .A(S), .Y(SB) );
  ND2_1959 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1958 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1957 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_652 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_652 UIV ( .A(S), .Y(SB) );
  ND2_1956 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1955 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1954 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_651 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_651 UIV ( .A(S), .Y(SB) );
  ND2_1953 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1952 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1951 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_650 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_650 UIV ( .A(S), .Y(SB) );
  ND2_1950 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1949 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1948 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_649 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_649 UIV ( .A(S), .Y(SB) );
  ND2_1947 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1946 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1945 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_648 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_648 UIV ( .A(S), .Y(SB) );
  ND2_1944 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1943 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1942 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_645 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_645 UIV ( .A(S), .Y(SB) );
  ND2_1935 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1934 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1933 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_641 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_641 UIV ( .A(S), .Y(SB) );
  ND2_1923 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1922 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1921 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_639 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_639 UIV ( .A(S), .Y(SB) );
  ND2_1917 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1916 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1915 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_637 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_637 UIV ( .A(S), .Y(SB) );
  ND2_1911 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1910 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1909 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_635 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_635 UIV ( .A(S), .Y(SB) );
  ND2_1905 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1904 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1903 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_633 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_633 UIV ( .A(S), .Y(SB) );
  ND2_1899 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1898 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1897 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_632 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_632 UIV ( .A(S), .Y(SB) );
  ND2_1896 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1895 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1894 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_631 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_631 UIV ( .A(S), .Y(SB) );
  ND2_1893 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1892 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1891 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_630 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_630 UIV ( .A(S), .Y(SB) );
  ND2_1890 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1889 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1888 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_629 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_629 UIV ( .A(S), .Y(SB) );
  ND2_1887 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1886 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1885 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_628 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_628 UIV ( .A(S), .Y(SB) );
  ND2_1884 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1883 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1882 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_627 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_627 UIV ( .A(S), .Y(SB) );
  ND2_1881 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1880 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1879 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_626 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_626 UIV ( .A(S), .Y(SB) );
  ND2_1878 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1877 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1876 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_625 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_625 UIV ( .A(S), .Y(SB) );
  ND2_1875 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1874 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1873 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_624 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_624 UIV ( .A(S), .Y(SB) );
  ND2_1872 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1871 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1870 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_623 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_623 UIV ( .A(S), .Y(SB) );
  ND2_1869 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1868 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1867 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_622 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_622 UIV ( .A(S), .Y(SB) );
  ND2_1866 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1865 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1864 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_621 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_621 UIV ( .A(S), .Y(SB) );
  ND2_1863 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1862 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1861 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_620 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_620 UIV ( .A(S), .Y(SB) );
  ND2_1860 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1859 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1858 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_619 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_619 UIV ( .A(S), .Y(SB) );
  ND2_1857 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1856 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1855 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_618 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_618 UIV ( .A(S), .Y(SB) );
  ND2_1854 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1853 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1852 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_617 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_617 UIV ( .A(S), .Y(SB) );
  ND2_1851 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1850 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1849 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_616 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_616 UIV ( .A(S), .Y(SB) );
  ND2_1848 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1847 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1846 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_615 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_615 UIV ( .A(S), .Y(SB) );
  ND2_1845 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1844 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1843 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_614 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_614 UIV ( .A(S), .Y(SB) );
  ND2_1842 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1841 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1840 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_613 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_613 UIV ( .A(S), .Y(SB) );
  ND2_1839 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1838 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1837 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_612 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_612 UIV ( .A(S), .Y(SB) );
  ND2_1836 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1835 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1834 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_611 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_611 UIV ( .A(S), .Y(SB) );
  ND2_1833 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1832 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1831 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_610 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_610 UIV ( .A(S), .Y(SB) );
  ND2_1830 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1829 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1828 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_609 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_609 UIV ( .A(S), .Y(SB) );
  ND2_1827 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1826 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1825 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_608 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_608 UIV ( .A(S), .Y(SB) );
  ND2_1824 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1823 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1822 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_607 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_607 UIV ( .A(S), .Y(SB) );
  ND2_1821 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1820 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1819 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_606 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_606 UIV ( .A(S), .Y(SB) );
  ND2_1818 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1817 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1816 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_605 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_605 UIV ( .A(S), .Y(SB) );
  ND2_1815 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1814 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1813 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_604 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_604 UIV ( .A(S), .Y(SB) );
  ND2_1812 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1811 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1810 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_603 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_603 UIV ( .A(S), .Y(SB) );
  ND2_1809 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1808 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1807 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_602 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_602 UIV ( .A(S), .Y(SB) );
  ND2_1806 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1805 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1804 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_601 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_601 UIV ( .A(S), .Y(SB) );
  ND2_1803 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1802 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1801 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_600 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_600 UIV ( .A(S), .Y(SB) );
  ND2_1800 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1799 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1798 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_599 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_599 UIV ( .A(S), .Y(SB) );
  ND2_1797 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1796 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1795 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_598 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_598 UIV ( .A(S), .Y(SB) );
  ND2_1794 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1793 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1792 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_597 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_597 UIV ( .A(S), .Y(SB) );
  ND2_1791 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1790 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1789 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_596 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_596 UIV ( .A(S), .Y(SB) );
  ND2_1788 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1787 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1786 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_595 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_595 UIV ( .A(S), .Y(SB) );
  ND2_1785 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1784 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1783 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_594 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_594 UIV ( .A(S), .Y(SB) );
  ND2_1782 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1781 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1780 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_593 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_593 UIV ( .A(S), .Y(SB) );
  ND2_1779 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1778 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1777 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_592 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_592 UIV ( .A(S), .Y(SB) );
  ND2_1776 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1775 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1774 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_591 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_591 UIV ( .A(S), .Y(SB) );
  ND2_1773 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1772 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1771 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_590 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_590 UIV ( .A(S), .Y(SB) );
  ND2_1770 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1769 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1768 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_589 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_589 UIV ( .A(S), .Y(SB) );
  ND2_1767 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1766 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1765 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_588 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_588 UIV ( .A(S), .Y(SB) );
  ND2_1764 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1763 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1762 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_587 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_587 UIV ( .A(S), .Y(SB) );
  ND2_1761 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1760 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1759 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_586 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_586 UIV ( .A(S), .Y(SB) );
  ND2_1758 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1757 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1756 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_585 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_585 UIV ( .A(S), .Y(SB) );
  ND2_1755 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1754 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1753 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_584 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_584 UIV ( .A(S), .Y(SB) );
  ND2_1752 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1751 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1750 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_583 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_583 UIV ( .A(S), .Y(SB) );
  ND2_1749 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1748 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1747 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_582 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_582 UIV ( .A(S), .Y(SB) );
  ND2_1746 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1745 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1744 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_581 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_581 UIV ( .A(S), .Y(SB) );
  ND2_1743 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1742 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1741 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_580 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_580 UIV ( .A(S), .Y(SB) );
  ND2_1740 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1739 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1738 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_579 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_579 UIV ( .A(S), .Y(SB) );
  ND2_1737 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1736 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1735 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_578 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_578 UIV ( .A(S), .Y(SB) );
  ND2_1734 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1733 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1732 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_577 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_577 UIV ( .A(S), .Y(SB) );
  ND2_1731 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1730 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1729 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_480 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_480 UIV ( .A(S), .Y(SB) );
  ND2_1440 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1439 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1438 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_479 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_479 UIV ( .A(S), .Y(SB) );
  ND2_1437 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1436 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1435 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_478 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_478 UIV ( .A(S), .Y(SB) );
  ND2_1434 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1433 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1432 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_477 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_477 UIV ( .A(S), .Y(SB) );
  ND2_1431 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1430 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1429 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_476 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_476 UIV ( .A(S), .Y(SB) );
  ND2_1428 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1427 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1426 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_475 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_475 UIV ( .A(S), .Y(SB) );
  ND2_1425 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1424 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1423 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_474 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_474 UIV ( .A(S), .Y(SB) );
  ND2_1422 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1421 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1420 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_473 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_473 UIV ( .A(S), .Y(SB) );
  ND2_1419 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1418 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1417 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_472 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_472 UIV ( .A(S), .Y(SB) );
  ND2_1416 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1415 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1414 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_471 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_471 UIV ( .A(S), .Y(SB) );
  ND2_1413 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1412 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1411 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_470 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_470 UIV ( .A(S), .Y(SB) );
  ND2_1410 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1409 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1408 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_469 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_469 UIV ( .A(S), .Y(SB) );
  ND2_1407 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1406 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1405 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_468 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_468 UIV ( .A(S), .Y(SB) );
  ND2_1404 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1403 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1402 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_467 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_467 UIV ( .A(S), .Y(SB) );
  ND2_1401 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1400 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1399 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_466 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_466 UIV ( .A(S), .Y(SB) );
  ND2_1398 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1397 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1396 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_465 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_465 UIV ( .A(S), .Y(SB) );
  ND2_1395 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1394 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1393 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_464 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_464 UIV ( .A(S), .Y(SB) );
  ND2_1392 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1391 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1390 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_463 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_463 UIV ( .A(S), .Y(SB) );
  ND2_1389 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1388 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1387 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_462 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_462 UIV ( .A(S), .Y(SB) );
  ND2_1386 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1385 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1384 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_461 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_461 UIV ( .A(S), .Y(SB) );
  ND2_1383 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1382 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1381 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_460 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_460 UIV ( .A(S), .Y(SB) );
  ND2_1380 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1379 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1378 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_459 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_459 UIV ( .A(S), .Y(SB) );
  ND2_1377 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1376 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1375 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_458 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_458 UIV ( .A(S), .Y(SB) );
  ND2_1374 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1373 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1372 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_457 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_457 UIV ( .A(S), .Y(SB) );
  ND2_1371 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1370 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1369 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_456 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_456 UIV ( .A(S), .Y(SB) );
  ND2_1368 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1367 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1366 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_455 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_455 UIV ( .A(S), .Y(SB) );
  ND2_1365 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1364 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1363 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_454 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_454 UIV ( .A(S), .Y(SB) );
  ND2_1362 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1361 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1360 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_453 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_453 UIV ( .A(S), .Y(SB) );
  ND2_1359 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1358 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1357 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_452 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_452 UIV ( .A(S), .Y(SB) );
  ND2_1356 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1355 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1354 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_451 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_451 UIV ( .A(S), .Y(SB) );
  ND2_1353 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1352 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1351 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_450 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_450 UIV ( .A(S), .Y(SB) );
  ND2_1350 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1349 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1348 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_449 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_449 UIV ( .A(S), .Y(SB) );
  ND2_1347 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1346 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1345 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_448 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_448 UIV ( .A(S), .Y(SB) );
  ND2_1344 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1343 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1342 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_447 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_447 UIV ( .A(S), .Y(SB) );
  ND2_1341 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1340 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1339 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_446 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_446 UIV ( .A(S), .Y(SB) );
  ND2_1338 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1337 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1336 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_445 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_445 UIV ( .A(S), .Y(SB) );
  ND2_1335 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1334 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1333 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_444 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_444 UIV ( .A(S), .Y(SB) );
  ND2_1332 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1331 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1330 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_443 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_443 UIV ( .A(S), .Y(SB) );
  ND2_1329 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1328 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1327 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_442 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_442 UIV ( .A(S), .Y(SB) );
  ND2_1326 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1325 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1324 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_441 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_441 UIV ( .A(S), .Y(SB) );
  ND2_1323 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1322 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1321 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_440 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_440 UIV ( .A(S), .Y(SB) );
  ND2_1320 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1319 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1318 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_439 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_439 UIV ( .A(S), .Y(SB) );
  ND2_1317 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1316 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1315 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_438 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_438 UIV ( .A(S), .Y(SB) );
  ND2_1314 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1313 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1312 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_437 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_437 UIV ( .A(S), .Y(SB) );
  ND2_1311 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1310 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1309 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_436 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_436 UIV ( .A(S), .Y(SB) );
  ND2_1308 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1307 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1306 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_435 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_435 UIV ( .A(S), .Y(SB) );
  ND2_1305 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1304 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1303 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_434 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_434 UIV ( .A(S), .Y(SB) );
  ND2_1302 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1301 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1300 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_433 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_433 UIV ( .A(S), .Y(SB) );
  ND2_1299 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1298 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1297 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_432 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_432 UIV ( .A(S), .Y(SB) );
  ND2_1296 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1295 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1294 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_431 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_431 UIV ( .A(S), .Y(SB) );
  ND2_1293 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1292 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1291 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_430 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_430 UIV ( .A(S), .Y(SB) );
  ND2_1290 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1289 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1288 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_429 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_429 UIV ( .A(S), .Y(SB) );
  ND2_1287 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1286 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1285 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_428 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_428 UIV ( .A(S), .Y(SB) );
  ND2_1284 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1283 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1282 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_427 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_427 UIV ( .A(S), .Y(SB) );
  ND2_1281 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1280 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1279 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_426 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_426 UIV ( .A(S), .Y(SB) );
  ND2_1278 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1277 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1276 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_425 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_425 UIV ( .A(S), .Y(SB) );
  ND2_1275 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1274 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1273 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_424 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_424 UIV ( .A(S), .Y(SB) );
  ND2_1272 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1271 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1270 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_423 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_423 UIV ( .A(S), .Y(SB) );
  ND2_1269 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1268 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1267 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_422 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_422 UIV ( .A(S), .Y(SB) );
  ND2_1266 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1265 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1264 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_421 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_421 UIV ( .A(S), .Y(SB) );
  ND2_1263 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1262 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1261 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_420 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_420 UIV ( .A(S), .Y(SB) );
  ND2_1260 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1259 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1258 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_419 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_419 UIV ( .A(S), .Y(SB) );
  ND2_1257 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1256 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1255 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_418 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_418 UIV ( .A(S), .Y(SB) );
  ND2_1254 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1253 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1252 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_417 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_417 UIV ( .A(S), .Y(SB) );
  ND2_1251 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1250 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1249 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_416 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_416 UIV ( .A(S), .Y(SB) );
  ND2_1248 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1247 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1246 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_415 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_415 UIV ( .A(S), .Y(SB) );
  ND2_1245 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1244 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1243 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_414 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_414 UIV ( .A(S), .Y(SB) );
  ND2_1242 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1241 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1240 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_413 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_413 UIV ( .A(S), .Y(SB) );
  ND2_1239 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1238 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1237 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_412 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_412 UIV ( .A(S), .Y(SB) );
  ND2_1236 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1235 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1234 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_411 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_411 UIV ( .A(S), .Y(SB) );
  ND2_1233 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1232 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1231 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_410 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_410 UIV ( .A(S), .Y(SB) );
  ND2_1230 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1229 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1228 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_409 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_409 UIV ( .A(S), .Y(SB) );
  ND2_1227 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1226 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1225 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_408 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_408 UIV ( .A(S), .Y(SB) );
  ND2_1224 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1223 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1222 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_407 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_407 UIV ( .A(S), .Y(SB) );
  ND2_1221 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1220 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1219 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_406 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_406 UIV ( .A(S), .Y(SB) );
  ND2_1218 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1217 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1216 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_405 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_405 UIV ( .A(S), .Y(SB) );
  ND2_1215 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1214 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1213 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_404 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_404 UIV ( .A(S), .Y(SB) );
  ND2_1212 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1211 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1210 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_403 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_403 UIV ( .A(S), .Y(SB) );
  ND2_1209 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1208 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1207 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_402 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_402 UIV ( .A(S), .Y(SB) );
  ND2_1206 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1205 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1204 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_401 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_401 UIV ( .A(S), .Y(SB) );
  ND2_1203 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1202 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1201 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_400 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_400 UIV ( .A(S), .Y(SB) );
  ND2_1200 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1199 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1198 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_399 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_399 UIV ( .A(S), .Y(SB) );
  ND2_1197 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1196 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1195 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_398 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_398 UIV ( .A(S), .Y(SB) );
  ND2_1194 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1193 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1192 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_397 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_397 UIV ( .A(S), .Y(SB) );
  ND2_1191 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1190 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1189 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_396 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_396 UIV ( .A(S), .Y(SB) );
  ND2_1188 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1187 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1186 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_395 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_395 UIV ( .A(S), .Y(SB) );
  ND2_1185 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1184 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1183 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_394 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_394 UIV ( .A(S), .Y(SB) );
  ND2_1182 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1181 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1180 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_393 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_393 UIV ( .A(S), .Y(SB) );
  ND2_1179 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1178 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1177 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_392 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_392 UIV ( .A(S), .Y(SB) );
  ND2_1176 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1175 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1174 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_391 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_391 UIV ( .A(S), .Y(SB) );
  ND2_1173 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1172 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1171 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_390 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_390 UIV ( .A(S), .Y(SB) );
  ND2_1170 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1169 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1168 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_389 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_389 UIV ( .A(S), .Y(SB) );
  ND2_1167 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1166 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1165 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_388 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_388 UIV ( .A(S), .Y(SB) );
  ND2_1164 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1163 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1162 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_387 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_387 UIV ( .A(S), .Y(SB) );
  ND2_1161 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1160 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1159 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_386 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_386 UIV ( .A(S), .Y(SB) );
  ND2_1158 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1157 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1156 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_385 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_385 UIV ( .A(S), .Y(SB) );
  ND2_1155 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1154 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1153 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_384 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_384 UIV ( .A(S), .Y(SB) );
  ND2_1152 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1151 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1150 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_383 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_383 UIV ( .A(S), .Y(SB) );
  ND2_1149 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1148 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1147 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_382 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_382 UIV ( .A(S), .Y(SB) );
  ND2_1146 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1145 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1144 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_381 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_381 UIV ( .A(S), .Y(SB) );
  ND2_1143 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1142 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1141 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_380 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_380 UIV ( .A(S), .Y(SB) );
  ND2_1140 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1139 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1138 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_379 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_379 UIV ( .A(S), .Y(SB) );
  ND2_1137 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1136 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1135 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_378 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_378 UIV ( .A(S), .Y(SB) );
  ND2_1134 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1133 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1132 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_377 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_377 UIV ( .A(S), .Y(SB) );
  ND2_1131 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1130 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1129 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_376 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_376 UIV ( .A(S), .Y(SB) );
  ND2_1128 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1127 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1126 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_375 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_375 UIV ( .A(S), .Y(SB) );
  ND2_1125 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1124 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1123 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_374 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_374 UIV ( .A(S), .Y(SB) );
  ND2_1122 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1121 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1120 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_373 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_373 UIV ( .A(S), .Y(SB) );
  ND2_1119 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1118 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1117 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_372 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_372 UIV ( .A(S), .Y(SB) );
  ND2_1116 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1115 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1114 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_371 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_371 UIV ( .A(S), .Y(SB) );
  ND2_1113 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1112 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1111 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_370 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_370 UIV ( .A(S), .Y(SB) );
  ND2_1110 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1109 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1108 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_369 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_369 UIV ( .A(S), .Y(SB) );
  ND2_1107 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1106 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1105 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_368 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_368 UIV ( .A(S), .Y(SB) );
  ND2_1104 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1103 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1102 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_367 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_367 UIV ( .A(S), .Y(SB) );
  ND2_1101 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1100 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1099 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_366 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_366 UIV ( .A(S), .Y(SB) );
  ND2_1098 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1097 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1096 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_365 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_365 UIV ( .A(S), .Y(SB) );
  ND2_1095 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1094 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1093 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_364 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_364 UIV ( .A(S), .Y(SB) );
  ND2_1092 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1091 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1090 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_363 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_363 UIV ( .A(S), .Y(SB) );
  ND2_1089 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1088 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1087 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_362 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_362 UIV ( .A(S), .Y(SB) );
  ND2_1086 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1085 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1084 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_361 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_361 UIV ( .A(S), .Y(SB) );
  ND2_1083 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1082 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1081 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_360 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_360 UIV ( .A(S), .Y(SB) );
  ND2_1080 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1079 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1078 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_359 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_359 UIV ( .A(S), .Y(SB) );
  ND2_1077 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1076 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1075 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_358 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_358 UIV ( .A(S), .Y(SB) );
  ND2_1074 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1073 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1072 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_357 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_357 UIV ( .A(S), .Y(SB) );
  ND2_1071 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1070 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1069 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_356 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_356 UIV ( .A(S), .Y(SB) );
  ND2_1068 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1067 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1066 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_355 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_355 UIV ( .A(S), .Y(SB) );
  ND2_1065 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1064 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1063 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_354 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_354 UIV ( .A(S), .Y(SB) );
  ND2_1062 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1061 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1060 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_353 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_353 UIV ( .A(S), .Y(SB) );
  ND2_1059 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1058 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1057 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_352 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_352 UIV ( .A(S), .Y(SB) );
  ND2_1056 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1055 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1054 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_351 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_351 UIV ( .A(S), .Y(SB) );
  ND2_1053 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1052 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1051 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_350 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_350 UIV ( .A(S), .Y(SB) );
  ND2_1050 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1049 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1048 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_349 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_349 UIV ( .A(S), .Y(SB) );
  ND2_1047 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1046 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1045 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_348 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_348 UIV ( .A(S), .Y(SB) );
  ND2_1044 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1043 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1042 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_347 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_347 UIV ( .A(S), .Y(SB) );
  ND2_1041 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1040 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1039 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_346 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_346 UIV ( .A(S), .Y(SB) );
  ND2_1038 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1037 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1036 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_345 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_345 UIV ( .A(S), .Y(SB) );
  ND2_1035 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1034 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1033 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_344 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_344 UIV ( .A(S), .Y(SB) );
  ND2_1032 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1031 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1030 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_343 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_343 UIV ( .A(S), .Y(SB) );
  ND2_1029 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1028 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1027 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_342 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_342 UIV ( .A(S), .Y(SB) );
  ND2_1026 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1025 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1024 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_341 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_341 UIV ( .A(S), .Y(SB) );
  ND2_1023 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1022 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1021 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_340 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_340 UIV ( .A(S), .Y(SB) );
  ND2_1020 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1019 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1018 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_339 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_339 UIV ( .A(S), .Y(SB) );
  ND2_1017 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1016 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1015 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_338 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_338 UIV ( .A(S), .Y(SB) );
  ND2_1014 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1013 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1012 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_337 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_337 UIV ( .A(S), .Y(SB) );
  ND2_1011 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1010 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1009 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_336 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_336 UIV ( .A(S), .Y(SB) );
  ND2_1008 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1007 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1006 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_335 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_335 UIV ( .A(S), .Y(SB) );
  ND2_1005 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1004 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1003 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_334 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_334 UIV ( .A(S), .Y(SB) );
  ND2_1002 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1001 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1000 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_333 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_333 UIV ( .A(S), .Y(SB) );
  ND2_999 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_998 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_997 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_332 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_332 UIV ( .A(S), .Y(SB) );
  ND2_996 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_995 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_994 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_331 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_331 UIV ( .A(S), .Y(SB) );
  ND2_993 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_992 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_991 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_330 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_330 UIV ( .A(S), .Y(SB) );
  ND2_990 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_989 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_988 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_329 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_329 UIV ( .A(S), .Y(SB) );
  ND2_987 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_986 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_985 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_328 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_328 UIV ( .A(S), .Y(SB) );
  ND2_984 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_983 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_982 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_327 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_327 UIV ( .A(S), .Y(SB) );
  ND2_981 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_980 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_979 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_326 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_326 UIV ( .A(S), .Y(SB) );
  ND2_978 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_977 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_976 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_325 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_325 UIV ( .A(S), .Y(SB) );
  ND2_975 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_974 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_973 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_324 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_324 UIV ( .A(S), .Y(SB) );
  ND2_972 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_971 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_970 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_323 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_323 UIV ( .A(S), .Y(SB) );
  ND2_969 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_968 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_967 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_322 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_322 UIV ( .A(S), .Y(SB) );
  ND2_966 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_965 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_964 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_321 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_321 UIV ( .A(S), .Y(SB) );
  ND2_963 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_962 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_961 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_320 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_320 UIV ( .A(S), .Y(SB) );
  ND2_960 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_959 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_958 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_319 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_319 UIV ( .A(S), .Y(SB) );
  ND2_957 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_956 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_955 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_318 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_318 UIV ( .A(S), .Y(SB) );
  ND2_954 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_953 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_952 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_317 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_317 UIV ( .A(S), .Y(SB) );
  ND2_951 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_950 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_949 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_316 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_316 UIV ( .A(S), .Y(SB) );
  ND2_948 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_947 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_946 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_315 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_315 UIV ( .A(S), .Y(SB) );
  ND2_945 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_944 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_943 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_314 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_314 UIV ( .A(S), .Y(SB) );
  ND2_942 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_941 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_940 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_313 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_313 UIV ( .A(S), .Y(SB) );
  ND2_939 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_938 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_937 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_311 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_311 UIV ( .A(S), .Y(SB) );
  ND2_933 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_932 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_931 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_308 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_308 UIV ( .A(S), .Y(SB) );
  ND2_924 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_923 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_922 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_307 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_307 UIV ( .A(S), .Y(SB) );
  ND2_921 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_920 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_919 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_300 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_300 UIV ( .A(S), .Y(SB) );
  ND2_900 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_899 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_898 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_299 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_299 UIV ( .A(S), .Y(SB) );
  ND2_897 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_896 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_895 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_298 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_298 UIV ( .A(S), .Y(SB) );
  ND2_894 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_893 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_892 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_297 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_297 UIV ( .A(S), .Y(SB) );
  ND2_891 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_890 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_889 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_295 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_295 UIV ( .A(S), .Y(SB) );
  ND2_885 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_884 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_883 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_288 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_288 UIV ( .A(S), .Y(SB) );
  ND2_864 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_863 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_862 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_287 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_287 UIV ( .A(S), .Y(SB) );
  ND2_861 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_860 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_859 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_286 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_286 UIV ( .A(S), .Y(SB) );
  ND2_858 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_857 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_856 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_285 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_285 UIV ( .A(S), .Y(SB) );
  ND2_855 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_854 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_853 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_284 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_284 UIV ( .A(S), .Y(SB) );
  ND2_852 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_851 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_850 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_283 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_283 UIV ( .A(S), .Y(SB) );
  ND2_849 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_848 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_847 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_282 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_282 UIV ( .A(S), .Y(SB) );
  ND2_846 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_845 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_844 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_281 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_281 UIV ( .A(S), .Y(SB) );
  ND2_843 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_842 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_841 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_275 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_275 UIV ( .A(S), .Y(SB) );
  ND2_825 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_824 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_823 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_272 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_272 UIV ( .A(S), .Y(SB) );
  ND2_816 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_815 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_814 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_271 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_271 UIV ( .A(S), .Y(SB) );
  ND2_813 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_812 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_811 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_270 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_270 UIV ( .A(S), .Y(SB) );
  ND2_810 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_809 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_808 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_267 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_267 UIV ( .A(S), .Y(SB) );
  ND2_801 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_800 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_799 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_266 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_266 UIV ( .A(S), .Y(SB) );
  ND2_798 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_797 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_796 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_265 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_265 UIV ( .A(S), .Y(SB) );
  ND2_795 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_794 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_793 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_264 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_264 UIV ( .A(S), .Y(SB) );
  ND2_792 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_791 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_790 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_263 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_263 UIV ( .A(S), .Y(SB) );
  ND2_789 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_788 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_787 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_256 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_256 UIV ( .A(S), .Y(SB) );
  ND2_768 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_767 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_766 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_255 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_255 UIV ( .A(S), .Y(SB) );
  ND2_765 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_764 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_763 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_254 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_254 UIV ( .A(S), .Y(SB) );
  ND2_762 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_761 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_760 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_253 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_253 UIV ( .A(S), .Y(SB) );
  ND2_759 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_758 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_757 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_252 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_252 UIV ( .A(S), .Y(SB) );
  ND2_756 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_755 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_754 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_251 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_251 UIV ( .A(S), .Y(SB) );
  ND2_753 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_752 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_751 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_250 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_250 UIV ( .A(S), .Y(SB) );
  ND2_750 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_749 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_748 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_249 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_249 UIV ( .A(S), .Y(SB) );
  ND2_747 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_746 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_745 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_248 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_248 UIV ( .A(S), .Y(SB) );
  ND2_744 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_743 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_742 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_247 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_247 UIV ( .A(S), .Y(SB) );
  ND2_741 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_740 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_739 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_246 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_246 UIV ( .A(S), .Y(SB) );
  ND2_738 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_737 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_736 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_245 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_245 UIV ( .A(S), .Y(SB) );
  ND2_735 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_734 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_733 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_244 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_244 UIV ( .A(S), .Y(SB) );
  ND2_732 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_731 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_730 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_243 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_243 UIV ( .A(S), .Y(SB) );
  ND2_729 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_728 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_727 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_242 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_242 UIV ( .A(S), .Y(SB) );
  ND2_726 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_725 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_724 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_241 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_241 UIV ( .A(S), .Y(SB) );
  ND2_723 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_722 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_721 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_240 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_240 UIV ( .A(S), .Y(SB) );
  ND2_720 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_719 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_718 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_239 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_239 UIV ( .A(S), .Y(SB) );
  ND2_717 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_716 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_715 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_238 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_238 UIV ( .A(S), .Y(SB) );
  ND2_714 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_713 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_712 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_237 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_237 UIV ( .A(S), .Y(SB) );
  ND2_711 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_710 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_709 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_236 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_236 UIV ( .A(S), .Y(SB) );
  ND2_708 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_707 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_706 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_235 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_235 UIV ( .A(S), .Y(SB) );
  ND2_705 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_704 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_703 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_234 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_234 UIV ( .A(S), .Y(SB) );
  ND2_702 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_701 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_700 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_233 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_233 UIV ( .A(S), .Y(SB) );
  ND2_699 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_698 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_697 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_232 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_232 UIV ( .A(S), .Y(SB) );
  ND2_696 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_695 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_694 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_231 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_231 UIV ( .A(S), .Y(SB) );
  ND2_693 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_692 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_691 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_230 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_230 UIV ( .A(S), .Y(SB) );
  ND2_690 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_689 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_688 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_229 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_229 UIV ( .A(S), .Y(SB) );
  ND2_687 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_686 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_685 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_228 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_228 UIV ( .A(S), .Y(SB) );
  ND2_684 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_683 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_682 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_227 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_227 UIV ( .A(S), .Y(SB) );
  ND2_681 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_680 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_679 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_226 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_226 UIV ( .A(S), .Y(SB) );
  ND2_678 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_677 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_676 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_225 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_225 UIV ( .A(S), .Y(SB) );
  ND2_675 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_674 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_673 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_219 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_219 UIV ( .A(S), .Y(SB) );
  ND2_657 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_656 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_655 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_217 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_217 UIV ( .A(S), .Y(SB) );
  ND2_651 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_650 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_649 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_215 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_215 UIV ( .A(S), .Y(SB) );
  ND2_645 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_644 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_643 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_214 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_214 UIV ( .A(S), .Y(SB) );
  ND2_642 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_641 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_640 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_213 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_213 UIV ( .A(S), .Y(SB) );
  ND2_639 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_638 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_637 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_206 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_206 UIV ( .A(S), .Y(SB) );
  ND2_618 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_617 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_616 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_202 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_202 UIV ( .A(S), .Y(SB) );
  ND2_606 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_605 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_604 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_200 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_200 UIV ( .A(S), .Y(SB) );
  ND2_600 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_599 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_598 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_199 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_199 UIV ( .A(S), .Y(SB) );
  ND2_597 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_596 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_595 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_198 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_198 UIV ( .A(S), .Y(SB) );
  ND2_594 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_593 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_592 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_197 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_197 UIV ( .A(S), .Y(SB) );
  ND2_591 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_590 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_589 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_196 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_196 UIV ( .A(S), .Y(SB) );
  ND2_588 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_587 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_586 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_195 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_195 UIV ( .A(S), .Y(SB) );
  ND2_585 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_584 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_583 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_194 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_194 UIV ( .A(S), .Y(SB) );
  ND2_582 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_581 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_580 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_193 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_193 UIV ( .A(S), .Y(SB) );
  ND2_579 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_578 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_577 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_192 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_192 UIV ( .A(S), .Y(SB) );
  ND2_576 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_575 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_574 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_189 UIV ( .A(S), .Y(SB) );
  ND2_567 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_566 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_565 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_187 UIV ( .A(S), .Y(SB) );
  ND2_561 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_560 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_559 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_186 UIV ( .A(S), .Y(SB) );
  ND2_558 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_557 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_556 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_183 UIV ( .A(S), .Y(SB) );
  ND2_549 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_548 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_547 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_177 UIV ( .A(S), .Y(SB) );
  ND2_531 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_530 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_529 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_174 UIV ( .A(S), .Y(SB) );
  ND2_522 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_521 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_520 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_169 UIV ( .A(S), .Y(SB) );
  ND2_507 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_506 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_505 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_167 UIV ( .A(S), .Y(SB) );
  ND2_501 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_500 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_499 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_166 UIV ( .A(S), .Y(SB) );
  ND2_498 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_497 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_496 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_165 UIV ( .A(S), .Y(SB) );
  ND2_495 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_494 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_493 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_164 UIV ( .A(S), .Y(SB) );
  ND2_492 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_491 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_490 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_163 UIV ( .A(S), .Y(SB) );
  ND2_489 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_488 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_487 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_162 UIV ( .A(S), .Y(SB) );
  ND2_486 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_485 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_484 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_161 UIV ( .A(S), .Y(SB) );
  ND2_483 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_482 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_481 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_160 UIV ( .A(S), .Y(SB) );
  ND2_480 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_479 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_478 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_158 UIV ( .A(S), .Y(SB) );
  ND2_474 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_473 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_472 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_155 UIV ( .A(S), .Y(SB) );
  ND2_465 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_464 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_463 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_153 UIV ( .A(S), .Y(SB) );
  ND2_459 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_458 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_457 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_151 UIV ( .A(S), .Y(SB) );
  ND2_453 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_452 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_451 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_150 UIV ( .A(S), .Y(SB) );
  ND2_450 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_449 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_448 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_149 UIV ( .A(S), .Y(SB) );
  ND2_447 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_446 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_445 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_142 UIV ( .A(S), .Y(SB) );
  ND2_426 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_425 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_424 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_137 UIV ( .A(S), .Y(SB) );
  ND2_411 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_410 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_409 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_134 UIV ( .A(S), .Y(SB) );
  ND2_402 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_401 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_400 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_133 UIV ( .A(S), .Y(SB) );
  ND2_399 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_398 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_397 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_132 UIV ( .A(S), .Y(SB) );
  ND2_396 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_395 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_394 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_131 UIV ( .A(S), .Y(SB) );
  ND2_393 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_392 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_391 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_130 UIV ( .A(S), .Y(SB) );
  ND2_390 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_389 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_388 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_129 UIV ( .A(S), .Y(SB) );
  ND2_387 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_386 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_385 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_128 UIV ( .A(S), .Y(SB) );
  ND2_384 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_383 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_382 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_127 UIV ( .A(S), .Y(SB) );
  ND2_381 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_380 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_379 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_126 UIV ( .A(S), .Y(SB) );
  ND2_378 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_377 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_376 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_123 UIV ( .A(S), .Y(SB) );
  ND2_369 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_368 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_367 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_122 UIV ( .A(S), .Y(SB) );
  ND2_366 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_365 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_364 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_117 UIV ( .A(S), .Y(SB) );
  ND2_351 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_350 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_349 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_113 UIV ( .A(S), .Y(SB) );
  ND2_339 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_338 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_337 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_111 UIV ( .A(S), .Y(SB) );
  ND2_333 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_332 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_331 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_105 UIV ( .A(S), .Y(SB) );
  ND2_315 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_314 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_313 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_101 UIV ( .A(S), .Y(SB) );
  ND2_303 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_302 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_301 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_99 UIV ( .A(S), .Y(SB) );
  ND2_297 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_296 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_295 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_98 UIV ( .A(S), .Y(SB) );
  ND2_294 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_293 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_292 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_97 UIV ( .A(S), .Y(SB) );
  ND2_291 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_290 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_289 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_96 UIV ( .A(S), .Y(SB) );
  ND2_288 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_287 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_286 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_95 UIV ( .A(S), .Y(SB) );
  ND2_285 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_284 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_283 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_94 UIV ( .A(S), .Y(SB) );
  ND2_282 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_281 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_280 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_93 UIV ( .A(S), .Y(SB) );
  ND2_279 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_278 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_277 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_91 UIV ( .A(S), .Y(SB) );
  ND2_273 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_272 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_271 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_89 UIV ( .A(S), .Y(SB) );
  ND2_267 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_266 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_265 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_86 UIV ( .A(S), .Y(SB) );
  ND2_258 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_257 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_256 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_82 UIV ( .A(S), .Y(SB) );
  ND2_246 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_245 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_244 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_79 UIV ( .A(S), .Y(SB) );
  ND2_237 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_236 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_235 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_78 UIV ( .A(S), .Y(SB) );
  ND2_234 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_233 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_232 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_70 UIV ( .A(S), .Y(SB) );
  ND2_210 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_209 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_208 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_67 UIV ( .A(S), .Y(SB) );
  ND2_201 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_200 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_199 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_65 UIV ( .A(S), .Y(SB) );
  ND2_195 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_194 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_193 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_64 UIV ( .A(S), .Y(SB) );
  ND2_192 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_191 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_190 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_63 UIV ( .A(S), .Y(SB) );
  ND2_189 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_188 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_187 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_62 UIV ( .A(S), .Y(SB) );
  ND2_186 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_185 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_184 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_61 UIV ( .A(S), .Y(SB) );
  ND2_183 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_182 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_181 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_59 UIV ( .A(S), .Y(SB) );
  ND2_177 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_176 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_175 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_58 UIV ( .A(S), .Y(SB) );
  ND2_174 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_173 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_172 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_57 UIV ( .A(S), .Y(SB) );
  ND2_171 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_170 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_169 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_50 UIV ( .A(S), .Y(SB) );
  ND2_150 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_149 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_148 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_49 UIV ( .A(S), .Y(SB) );
  ND2_147 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_146 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_145 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_46 UIV ( .A(S), .Y(SB) );
  ND2_138 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_137 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_136 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_45 UIV ( .A(S), .Y(SB) );
  ND2_135 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_134 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_133 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_41 UIV ( .A(S), .Y(SB) );
  ND2_123 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_122 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_121 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_37 UIV ( .A(S), .Y(SB) );
  ND2_111 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_110 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_109 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_34 UIV ( .A(S), .Y(SB) );
  ND2_102 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_101 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_100 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_33 UIV ( .A(S), .Y(SB) );
  ND2_99 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_98 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_97 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_32 UIV ( .A(S), .Y(SB) );
  ND2_96 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_95 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_94 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_31 UIV ( .A(S), .Y(SB) );
  ND2_93 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_92 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_91 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_30 UIV ( .A(S), .Y(SB) );
  ND2_90 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_89 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_88 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_29 UIV ( .A(S), .Y(SB) );
  ND2_87 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_86 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_85 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_28 UIV ( .A(S), .Y(SB) );
  ND2_84 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_83 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_82 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_27 UIV ( .A(S), .Y(SB) );
  ND2_81 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_80 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_79 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_26 UIV ( .A(S), .Y(SB) );
  ND2_78 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_77 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_76 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_25 UIV ( .A(S), .Y(SB) );
  ND2_75 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_74 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_73 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_22 UIV ( .A(S), .Y(SB) );
  ND2_66 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_65 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_64 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_21 UIV ( .A(S), .Y(SB) );
  ND2_63 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_62 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_61 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_17 UIV ( .A(S), .Y(SB) );
  ND2_51 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_50 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_49 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_14 UIV ( .A(S), .Y(SB) );
  ND2_42 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_41 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_40 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_13 UIV ( .A(S), .Y(SB) );
  ND2_39 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_38 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_37 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_10 UIV ( .A(S), .Y(SB) );
  ND2_30 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_29 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_28 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_9 UIV ( .A(S), .Y(SB) );
  ND2_27 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_26 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_25 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_5 UIV ( .A(S), .Y(SB) );
  ND2_15 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_14 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_13 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_920 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_920 UIV ( .A(S), .Y(SB) );
  ND2_2760 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2759 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2758 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_735 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_735 UIV ( .A(S), .Y(SB) );
  ND2_2205 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2204 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2203 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_732 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_732 UIV ( .A(S), .Y(SB) );
  ND2_2196 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2195 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2194 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_711 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_711 UIV ( .A(S), .Y(SB) );
  ND2_2133 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2132 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2131 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_709 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_709 UIV ( .A(S), .Y(SB) );
  ND2_2127 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2126 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2125 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_312 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_312 UIV ( .A(S), .Y(SB) );
  ND2_936 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_935 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_934 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_310 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_310 UIV ( .A(S), .Y(SB) );
  ND2_930 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_929 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_928 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_309 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_309 UIV ( .A(S), .Y(SB) );
  ND2_927 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_926 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_925 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_306 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_306 UIV ( .A(S), .Y(SB) );
  ND2_918 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_917 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_916 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_305 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_305 UIV ( .A(S), .Y(SB) );
  ND2_915 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_914 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_913 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_304 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_304 UIV ( .A(S), .Y(SB) );
  ND2_912 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_911 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_910 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_303 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_303 UIV ( .A(S), .Y(SB) );
  ND2_909 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_908 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_907 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_302 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_302 UIV ( .A(S), .Y(SB) );
  ND2_906 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_905 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_904 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_301 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_301 UIV ( .A(S), .Y(SB) );
  ND2_903 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_902 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_901 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_296 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_296 UIV ( .A(S), .Y(SB) );
  ND2_888 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_887 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_886 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_294 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_294 UIV ( .A(S), .Y(SB) );
  ND2_882 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_881 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_880 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_293 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_293 UIV ( .A(S), .Y(SB) );
  ND2_879 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_878 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_877 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_292 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_292 UIV ( .A(S), .Y(SB) );
  ND2_876 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_875 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_874 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_291 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_291 UIV ( .A(S), .Y(SB) );
  ND2_873 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_872 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_871 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_290 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_290 UIV ( .A(S), .Y(SB) );
  ND2_870 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_869 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_868 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_289 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_289 UIV ( .A(S), .Y(SB) );
  ND2_867 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_866 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_865 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_280 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_280 UIV ( .A(S), .Y(SB) );
  ND2_840 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_839 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_838 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_279 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_279 UIV ( .A(S), .Y(SB) );
  ND2_837 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_836 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_835 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_278 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_278 UIV ( .A(S), .Y(SB) );
  ND2_834 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_833 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_832 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_277 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_277 UIV ( .A(S), .Y(SB) );
  ND2_831 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_830 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_829 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_276 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_276 UIV ( .A(S), .Y(SB) );
  ND2_828 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_827 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_826 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_274 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_274 UIV ( .A(S), .Y(SB) );
  ND2_822 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_821 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_820 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_273 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_273 UIV ( .A(S), .Y(SB) );
  ND2_819 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_818 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_817 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_269 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_269 UIV ( .A(S), .Y(SB) );
  ND2_807 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_806 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_805 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_268 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_268 UIV ( .A(S), .Y(SB) );
  ND2_804 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_803 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_802 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_262 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_262 UIV ( .A(S), .Y(SB) );
  ND2_786 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_785 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_784 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_261 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_261 UIV ( .A(S), .Y(SB) );
  ND2_783 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_782 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_781 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_260 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_260 UIV ( .A(S), .Y(SB) );
  ND2_780 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_779 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_778 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_259 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_259 UIV ( .A(S), .Y(SB) );
  ND2_777 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_776 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_775 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_258 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_258 UIV ( .A(S), .Y(SB) );
  ND2_774 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_773 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_772 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_257 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_257 UIV ( .A(S), .Y(SB) );
  ND2_771 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_770 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_769 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_224 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_224 UIV ( .A(S), .Y(SB) );
  ND2_672 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_671 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_670 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_222 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_222 UIV ( .A(S), .Y(SB) );
  ND2_666 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_665 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_664 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_221 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_221 UIV ( .A(S), .Y(SB) );
  ND2_663 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_662 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_661 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_201 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_201 UIV ( .A(S), .Y(SB) );
  ND2_603 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_602 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_601 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_185 UIV ( .A(S), .Y(SB) );
  ND2_555 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_554 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_553 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_181 UIV ( .A(S), .Y(SB) );
  ND2_543 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_542 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_541 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_145 UIV ( .A(S), .Y(SB) );
  ND2_435 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_434 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_433 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_141 UIV ( .A(S), .Y(SB) );
  ND2_423 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_422 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_421 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_121 UIV ( .A(S), .Y(SB) );
  ND2_363 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_362 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_361 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_85 UIV ( .A(S), .Y(SB) );
  ND2_255 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_254 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_253 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_73 UIV ( .A(S), .Y(SB) );
  ND2_219 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_218 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_217 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_69 UIV ( .A(S), .Y(SB) );
  ND2_207 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_206 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_205 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_741 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_741 UIV ( .A(S), .Y(SB) );
  ND2_2223 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2222 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2221 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_740 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_740 UIV ( .A(S), .Y(SB) );
  ND2_2220 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2219 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2218 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_739 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_739 UIV ( .A(S), .Y(SB) );
  ND2_2217 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2216 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2215 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_729 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_729 UIV ( .A(S), .Y(SB) );
  ND2_2187 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2186 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2185 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_725 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_725 UIV ( .A(S), .Y(SB) );
  ND2_2175 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2174 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2173 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_724 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_724 UIV ( .A(S), .Y(SB) );
  ND2_2172 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2171 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2170 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_715 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_715 UIV ( .A(S), .Y(SB) );
  ND2_2145 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2144 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2143 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_714 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_714 UIV ( .A(S), .Y(SB) );
  ND2_2142 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2141 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2140 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_713 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_713 UIV ( .A(S), .Y(SB) );
  ND2_2139 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2138 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2137 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_646 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_646 UIV ( .A(S), .Y(SB) );
  ND2_1938 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1937 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1936 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_644 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_644 UIV ( .A(S), .Y(SB) );
  ND2_1932 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1931 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1930 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_643 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_643 UIV ( .A(S), .Y(SB) );
  ND2_1929 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1928 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1927 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_642 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_642 UIV ( .A(S), .Y(SB) );
  ND2_1926 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1925 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1924 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_640 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_640 UIV ( .A(S), .Y(SB) );
  ND2_1920 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1919 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1918 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_638 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_638 UIV ( .A(S), .Y(SB) );
  ND2_1914 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1913 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1912 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_636 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_636 UIV ( .A(S), .Y(SB) );
  ND2_1908 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1907 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1906 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_634 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_634 UIV ( .A(S), .Y(SB) );
  ND2_1902 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1901 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1900 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_223 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_223 UIV ( .A(S), .Y(SB) );
  ND2_669 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_668 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_667 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_218 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_218 UIV ( .A(S), .Y(SB) );
  ND2_654 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_653 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_652 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_216 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_216 UIV ( .A(S), .Y(SB) );
  ND2_648 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_647 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_646 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_208 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_208 UIV ( .A(S), .Y(SB) );
  ND2_624 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_623 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_622 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_207 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_207 UIV ( .A(S), .Y(SB) );
  ND2_621 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_620 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_619 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_205 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_205 UIV ( .A(S), .Y(SB) );
  ND2_615 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_614 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_613 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_204 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_204 UIV ( .A(S), .Y(SB) );
  ND2_612 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_611 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_610 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_203 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_203 UIV ( .A(S), .Y(SB) );
  ND2_609 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_608 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_607 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_191 UIV ( .A(S), .Y(SB) );
  ND2_573 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_572 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_571 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_190 UIV ( .A(S), .Y(SB) );
  ND2_570 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_569 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_568 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_182 UIV ( .A(S), .Y(SB) );
  ND2_546 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_545 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_544 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_179 UIV ( .A(S), .Y(SB) );
  ND2_537 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_536 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_535 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_178 UIV ( .A(S), .Y(SB) );
  ND2_534 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_533 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_532 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_170 UIV ( .A(S), .Y(SB) );
  ND2_510 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_509 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_508 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_168 UIV ( .A(S), .Y(SB) );
  ND2_504 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_503 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_502 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_159 UIV ( .A(S), .Y(SB) );
  ND2_477 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_476 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_475 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_157 UIV ( .A(S), .Y(SB) );
  ND2_471 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_470 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_469 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_154 UIV ( .A(S), .Y(SB) );
  ND2_462 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_461 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_460 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_147 UIV ( .A(S), .Y(SB) );
  ND2_441 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_440 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_439 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_146 UIV ( .A(S), .Y(SB) );
  ND2_438 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_437 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_436 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_143 UIV ( .A(S), .Y(SB) );
  ND2_429 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_428 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_427 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_136 UIV ( .A(S), .Y(SB) );
  ND2_408 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_407 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_406 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_135 UIV ( .A(S), .Y(SB) );
  ND2_405 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_404 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_403 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_125 UIV ( .A(S), .Y(SB) );
  ND2_375 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_374 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_373 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_119 UIV ( .A(S), .Y(SB) );
  ND2_357 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_356 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_355 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_118 UIV ( .A(S), .Y(SB) );
  ND2_354 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_353 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_352 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_116 UIV ( .A(S), .Y(SB) );
  ND2_348 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_347 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_346 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_115 UIV ( .A(S), .Y(SB) );
  ND2_345 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_344 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_343 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_112 UIV ( .A(S), .Y(SB) );
  ND2_336 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_335 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_334 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_110 UIV ( .A(S), .Y(SB) );
  ND2_330 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_329 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_328 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_109 UIV ( .A(S), .Y(SB) );
  ND2_327 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_326 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_325 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_102 UIV ( .A(S), .Y(SB) );
  ND2_306 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_305 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_304 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_100 UIV ( .A(S), .Y(SB) );
  ND2_300 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_299 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_298 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_92 UIV ( .A(S), .Y(SB) );
  ND2_276 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_275 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_274 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_90 UIV ( .A(S), .Y(SB) );
  ND2_270 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_269 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_268 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_87 UIV ( .A(S), .Y(SB) );
  ND2_261 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_260 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_259 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_83 UIV ( .A(S), .Y(SB) );
  ND2_249 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_248 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_247 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_81 UIV ( .A(S), .Y(SB) );
  ND2_243 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_242 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_241 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_77 UIV ( .A(S), .Y(SB) );
  ND2_231 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_230 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_229 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_66 UIV ( .A(S), .Y(SB) );
  ND2_198 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_197 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_196 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_60 UIV ( .A(S), .Y(SB) );
  ND2_180 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_179 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_178 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_55 UIV ( .A(S), .Y(SB) );
  ND2_165 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_164 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_163 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_54 UIV ( .A(S), .Y(SB) );
  ND2_162 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_161 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_160 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_51 UIV ( .A(S), .Y(SB) );
  ND2_153 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_152 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_151 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_47 UIV ( .A(S), .Y(SB) );
  ND2_141 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_140 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_139 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_43 UIV ( .A(S), .Y(SB) );
  ND2_129 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_128 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_127 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_42 UIV ( .A(S), .Y(SB) );
  ND2_126 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_125 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_124 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_38 UIV ( .A(S), .Y(SB) );
  ND2_114 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_113 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_112 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_211 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_211 UIV ( .A(S), .Y(SB) );
  ND2_633 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_632 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_631 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_210 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_210 UIV ( .A(S), .Y(SB) );
  ND2_630 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_629 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_628 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_180 UIV ( .A(S), .Y(SB) );
  ND2_540 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_539 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_538 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_172 UIV ( .A(S), .Y(SB) );
  ND2_516 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_515 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_514 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_108 UIV ( .A(S), .Y(SB) );
  ND2_324 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_323 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_322 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_104 UIV ( .A(S), .Y(SB) );
  ND2_312 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_311 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_310 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_72 UIV ( .A(S), .Y(SB) );
  ND2_216 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_215 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_214 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_36 UIV ( .A(S), .Y(SB) );
  ND2_108 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_107 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_106 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_188 UIV ( .A(S), .Y(SB) );
  ND2_564 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_563 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_562 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_184 UIV ( .A(S), .Y(SB) );
  ND2_552 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_551 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_550 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_176 UIV ( .A(S), .Y(SB) );
  ND2_528 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_527 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_526 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_175 UIV ( .A(S), .Y(SB) );
  ND2_525 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_524 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_523 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_171 UIV ( .A(S), .Y(SB) );
  ND2_513 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_512 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_511 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_156 UIV ( .A(S), .Y(SB) );
  ND2_468 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_467 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_466 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_152 UIV ( .A(S), .Y(SB) );
  ND2_456 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_455 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_454 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_148 UIV ( .A(S), .Y(SB) );
  ND2_444 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_443 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_442 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_144 UIV ( .A(S), .Y(SB) );
  ND2_432 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_431 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_430 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_140 UIV ( .A(S), .Y(SB) );
  ND2_420 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_419 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_418 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_139 UIV ( .A(S), .Y(SB) );
  ND2_417 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_416 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_415 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_138 UIV ( .A(S), .Y(SB) );
  ND2_414 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_413 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_412 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_124 UIV ( .A(S), .Y(SB) );
  ND2_372 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_371 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_370 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_120 UIV ( .A(S), .Y(SB) );
  ND2_360 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_359 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_358 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_107 UIV ( .A(S), .Y(SB) );
  ND2_321 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_320 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_319 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_106 UIV ( .A(S), .Y(SB) );
  ND2_318 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_317 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_316 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_88 UIV ( .A(S), .Y(SB) );
  ND2_264 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_263 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_262 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_84 UIV ( .A(S), .Y(SB) );
  ND2_252 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_251 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_250 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_76 UIV ( .A(S), .Y(SB) );
  ND2_228 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_227 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_226 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_75 UIV ( .A(S), .Y(SB) );
  ND2_225 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_224 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_223 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_74 UIV ( .A(S), .Y(SB) );
  ND2_222 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_221 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_220 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_71 UIV ( .A(S), .Y(SB) );
  ND2_213 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_212 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_211 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_68 UIV ( .A(S), .Y(SB) );
  ND2_204 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_203 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_202 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_56 UIV ( .A(S), .Y(SB) );
  ND2_168 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_167 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_166 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_52 UIV ( .A(S), .Y(SB) );
  ND2_156 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_155 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_154 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_48 UIV ( .A(S), .Y(SB) );
  ND2_144 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_143 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_142 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_44 UIV ( .A(S), .Y(SB) );
  ND2_132 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_131 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_130 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_40 UIV ( .A(S), .Y(SB) );
  ND2_120 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_119 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_118 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_39 UIV ( .A(S), .Y(SB) );
  ND2_117 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_116 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_115 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_35 UIV ( .A(S), .Y(SB) );
  ND2_105 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_104 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_103 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_886 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_886 UIV ( .A(S), .Y(SB) );
  ND2_2658 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2657 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2656 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_885 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_885 UIV ( .A(S), .Y(SB) );
  ND2_2655 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2654 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2653 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_884 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_884 UIV ( .A(S), .Y(SB) );
  ND2_2652 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2651 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2650 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_883 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_883 UIV ( .A(S), .Y(SB) );
  ND2_2649 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2648 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2647 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_882 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_882 UIV ( .A(S), .Y(SB) );
  ND2_2646 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2645 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2644 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_881 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_881 UIV ( .A(S), .Y(SB) );
  ND2_2643 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2642 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2641 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_880 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_880 UIV ( .A(S), .Y(SB) );
  ND2_2640 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2639 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2638 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_879 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_879 UIV ( .A(S), .Y(SB) );
  ND2_2637 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2636 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2635 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_878 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_878 UIV ( .A(S), .Y(SB) );
  ND2_2634 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2633 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2632 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_877 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_877 UIV ( .A(S), .Y(SB) );
  ND2_2631 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2630 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2629 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_876 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_876 UIV ( .A(S), .Y(SB) );
  ND2_2628 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2627 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2626 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_875 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_875 UIV ( .A(S), .Y(SB) );
  ND2_2625 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2624 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2623 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_874 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_874 UIV ( .A(S), .Y(SB) );
  ND2_2622 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2621 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2620 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_873 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_873 UIV ( .A(S), .Y(SB) );
  ND2_2619 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2618 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2617 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_872 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_872 UIV ( .A(S), .Y(SB) );
  ND2_2616 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2615 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2614 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_871 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_871 UIV ( .A(S), .Y(SB) );
  ND2_2613 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2612 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2611 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_870 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_870 UIV ( .A(S), .Y(SB) );
  ND2_2610 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2609 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2608 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_869 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_869 UIV ( .A(S), .Y(SB) );
  ND2_2607 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2606 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2605 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_868 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_868 UIV ( .A(S), .Y(SB) );
  ND2_2604 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2603 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2602 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_867 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_867 UIV ( .A(S), .Y(SB) );
  ND2_2601 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2600 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2599 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_866 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_866 UIV ( .A(S), .Y(SB) );
  ND2_2598 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2597 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2596 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_865 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_865 UIV ( .A(S), .Y(SB) );
  ND2_2595 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2594 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2593 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_864 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_864 UIV ( .A(S), .Y(SB) );
  ND2_2592 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2591 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2590 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_863 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_863 UIV ( .A(S), .Y(SB) );
  ND2_2589 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2588 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2587 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_862 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_862 UIV ( .A(S), .Y(SB) );
  ND2_2586 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2585 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2584 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_861 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_861 UIV ( .A(S), .Y(SB) );
  ND2_2583 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2582 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2581 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_860 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_860 UIV ( .A(S), .Y(SB) );
  ND2_2580 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2579 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2578 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_859 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_859 UIV ( .A(S), .Y(SB) );
  ND2_2577 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2576 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2575 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_858 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_858 UIV ( .A(S), .Y(SB) );
  ND2_2574 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2573 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2572 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_857 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_857 UIV ( .A(S), .Y(SB) );
  ND2_2571 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2570 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2569 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_856 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_856 UIV ( .A(S), .Y(SB) );
  ND2_2568 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2567 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2566 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_806 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_806 UIV ( .A(S), .Y(SB) );
  ND2_2418 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2417 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2416 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_798 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_798 UIV ( .A(S), .Y(SB) );
  ND2_2394 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2393 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2392 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_770 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_770 UIV ( .A(S), .Y(SB) );
  ND2_2310 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2309 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2308 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_769 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_769 UIV ( .A(S), .Y(SB) );
  ND2_2307 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2306 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2305 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_209 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_209 UIV ( .A(S), .Y(SB) );
  ND2_627 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_626 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_625 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_173 UIV ( .A(S), .Y(SB) );
  ND2_519 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_518 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_517 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_114 UIV ( .A(S), .Y(SB) );
  ND2_342 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_341 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_340 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_103 UIV ( .A(S), .Y(SB) );
  ND2_309 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_308 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_307 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_24 UIV ( .A(S), .Y(SB) );
  ND2_72 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_71 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_70 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_23 UIV ( .A(S), .Y(SB) );
  ND2_69 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_68 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_67 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_20 UIV ( .A(S), .Y(SB) );
  ND2_60 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_59 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_58 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_19 UIV ( .A(S), .Y(SB) );
  ND2_57 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_56 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_55 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_18 UIV ( .A(S), .Y(SB) );
  ND2_54 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_53 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_52 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_16 UIV ( .A(S), .Y(SB) );
  ND2_48 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_47 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_46 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_12 UIV ( .A(S), .Y(SB) );
  ND2_36 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_35 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_34 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_11 UIV ( .A(S), .Y(SB) );
  ND2_33 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_32 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_31 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_8 UIV ( .A(S), .Y(SB) );
  ND2_24 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_23 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_22 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_7 UIV ( .A(S), .Y(SB) );
  ND2_21 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_20 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_19 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_6 UIV ( .A(S), .Y(SB) );
  ND2_18 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_17 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_16 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_4 UIV ( .A(S), .Y(SB) );
  ND2_12 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_11 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_10 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_3 UIV ( .A(S), .Y(SB) );
  ND2_9 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_8 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_7 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_2 UIV ( .A(S), .Y(SB) );
  ND2_6 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_5 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_4 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_1 UIV ( .A(S), .Y(SB) );
  ND2_3 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module D_Reg_generic_N32_6 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55837, net55838, net55839, net55840, net55841, net55842,
         net55843, net55844, net55845, net55846, net55847, net55848, net55849,
         net55850, net55851, net55852, net55853, net55854, net55855, net55856,
         net55857, net55858, net55859, net55860, net55861, net55862, net55863,
         net55864, net55865, net55866, net55867, net55868, n73, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146;
  assign n73 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n114), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n112), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n114), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n112), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n114), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n112), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n112), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n112), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n114), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n112), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n112), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n112), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n114), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n113), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n113), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n113), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n112), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n113), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n113), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n113), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n113), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n113), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n114), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n112), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n114), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n112), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n113), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n112), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n113), .Q(Q[3]), .QN(net55840)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n113), .Q(Q[2]), .QN(net55839)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n113), .Q(Q[1]), .QN(net55838)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n114), .Q(Q[0]), .QN(net55837)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n107) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n106) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n108) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n110) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n109) );
  OAI21_X1 U7 ( .B1(net55838), .B2(n108), .A(n139), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(n107), .ZN(n139) );
  OAI21_X1 U9 ( .B1(net55861), .B2(n108), .A(n145), .ZN(n8) );
  NAND2_X1 U10 ( .A1(D[24]), .A2(n106), .ZN(n145) );
  OAI21_X1 U11 ( .B1(net55862), .B2(n108), .A(n144), .ZN(n7) );
  NAND2_X1 U12 ( .A1(D[25]), .A2(n106), .ZN(n144) );
  OAI21_X1 U13 ( .B1(net55864), .B2(n108), .A(n142), .ZN(n5) );
  NAND2_X1 U14 ( .A1(D[27]), .A2(n106), .ZN(n142) );
  OAI21_X1 U15 ( .B1(net55865), .B2(n108), .A(n141), .ZN(n4) );
  NAND2_X1 U16 ( .A1(D[28]), .A2(n107), .ZN(n141) );
  OAI21_X1 U17 ( .B1(net55837), .B2(n109), .A(n140), .ZN(n32) );
  NAND2_X1 U18 ( .A1(D[0]), .A2(n107), .ZN(n140) );
  OAI21_X1 U19 ( .B1(net55839), .B2(n109), .A(n138), .ZN(n30) );
  NAND2_X1 U20 ( .A1(D[2]), .A2(n107), .ZN(n138) );
  OAI21_X1 U21 ( .B1(net55840), .B2(n109), .A(n136), .ZN(n29) );
  NAND2_X1 U22 ( .A1(D[3]), .A2(n107), .ZN(n136) );
  OAI21_X1 U23 ( .B1(net55847), .B2(n110), .A(n129), .ZN(n22) );
  NAND2_X1 U24 ( .A1(D[10]), .A2(n107), .ZN(n129) );
  OAI21_X1 U25 ( .B1(net55848), .B2(n110), .A(n128), .ZN(n21) );
  NAND2_X1 U26 ( .A1(D[11]), .A2(n107), .ZN(n128) );
  OAI21_X1 U27 ( .B1(net55849), .B2(n110), .A(n127), .ZN(n20) );
  NAND2_X1 U28 ( .A1(D[12]), .A2(n107), .ZN(n127) );
  OAI21_X1 U29 ( .B1(net55850), .B2(n110), .A(n125), .ZN(n19) );
  NAND2_X1 U30 ( .A1(D[13]), .A2(n107), .ZN(n125) );
  OAI21_X1 U31 ( .B1(net55851), .B2(n110), .A(n124), .ZN(n18) );
  NAND2_X1 U32 ( .A1(D[14]), .A2(n107), .ZN(n124) );
  OAI21_X1 U33 ( .B1(net55852), .B2(n110), .A(n123), .ZN(n17) );
  NAND2_X1 U34 ( .A1(D[15]), .A2(n107), .ZN(n123) );
  OAI21_X1 U35 ( .B1(net55853), .B2(n110), .A(n122), .ZN(n16) );
  NAND2_X1 U36 ( .A1(D[16]), .A2(n106), .ZN(n122) );
  OAI21_X1 U37 ( .B1(net55854), .B2(n110), .A(n121), .ZN(n15) );
  NAND2_X1 U38 ( .A1(D[17]), .A2(n106), .ZN(n121) );
  OAI21_X1 U39 ( .B1(net55855), .B2(n110), .A(n120), .ZN(n14) );
  NAND2_X1 U40 ( .A1(D[18]), .A2(n106), .ZN(n120) );
  OAI21_X1 U41 ( .B1(net55856), .B2(n110), .A(n119), .ZN(n13) );
  NAND2_X1 U42 ( .A1(D[19]), .A2(n106), .ZN(n119) );
  OAI21_X1 U43 ( .B1(net55863), .B2(n109), .A(n143), .ZN(n6) );
  NAND2_X1 U44 ( .A1(D[26]), .A2(n106), .ZN(n143) );
  OAI21_X1 U45 ( .B1(net55867), .B2(n110), .A(n126), .ZN(n2) );
  NAND2_X1 U46 ( .A1(D[30]), .A2(n107), .ZN(n126) );
  OAI21_X1 U47 ( .B1(net55868), .B2(n109), .A(n115), .ZN(n1) );
  NAND2_X1 U48 ( .A1(D[31]), .A2(n106), .ZN(n115) );
  OAI21_X1 U49 ( .B1(net55857), .B2(n111), .A(n118), .ZN(n12) );
  NAND2_X1 U50 ( .A1(D[20]), .A2(n106), .ZN(n118) );
  OAI21_X1 U51 ( .B1(net55858), .B2(n111), .A(n117), .ZN(n11) );
  NAND2_X1 U52 ( .A1(D[21]), .A2(n106), .ZN(n117) );
  OAI21_X1 U53 ( .B1(net55859), .B2(n111), .A(n116), .ZN(n10) );
  NAND2_X1 U54 ( .A1(D[22]), .A2(n106), .ZN(n116) );
  OAI21_X1 U55 ( .B1(net55841), .B2(n109), .A(n135), .ZN(n28) );
  NAND2_X1 U56 ( .A1(D[4]), .A2(n108), .ZN(n135) );
  OAI21_X1 U57 ( .B1(net55842), .B2(n109), .A(n134), .ZN(n27) );
  NAND2_X1 U58 ( .A1(D[5]), .A2(n108), .ZN(n134) );
  OAI21_X1 U59 ( .B1(net55843), .B2(n109), .A(n133), .ZN(n26) );
  NAND2_X1 U60 ( .A1(D[6]), .A2(n108), .ZN(n133) );
  OAI21_X1 U61 ( .B1(net55844), .B2(n109), .A(n132), .ZN(n25) );
  NAND2_X1 U62 ( .A1(D[7]), .A2(n108), .ZN(n132) );
  OAI21_X1 U63 ( .B1(net55845), .B2(n109), .A(n131), .ZN(n24) );
  NAND2_X1 U64 ( .A1(D[8]), .A2(n108), .ZN(n131) );
  OAI21_X1 U65 ( .B1(net55846), .B2(n110), .A(n130), .ZN(n23) );
  NAND2_X1 U66 ( .A1(D[9]), .A2(n108), .ZN(n130) );
  OAI21_X1 U67 ( .B1(net55866), .B2(n109), .A(n137), .ZN(n3) );
  NAND2_X1 U68 ( .A1(D[29]), .A2(n108), .ZN(n137) );
  OAI21_X1 U69 ( .B1(net55860), .B2(n109), .A(n146), .ZN(n9) );
  NAND2_X1 U70 ( .A1(n111), .A2(D[23]), .ZN(n146) );
  BUF_X1 U71 ( .A(n73), .Z(n113) );
  BUF_X1 U72 ( .A(n73), .Z(n112) );
  BUF_X1 U73 ( .A(n73), .Z(n114) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n111) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net179233, net232967, net243676, n10, n11, n12;
  assign Co = net179233;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n10) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n10), .ZN(n12) );
  NAND2_X1 U3 ( .A1(n12), .A2(n11), .ZN(net179233) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(net232967) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n11) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(net243676) );
  XNOR2_X1 U7 ( .A(net243676), .B(net232967), .ZN(S) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net179236, net240355, net241881, net223706, net223704, n8, n9, n10;
  assign Co = net179236;

  NAND2_X1 U1 ( .A1(net223706), .A2(Ci), .ZN(n9) );
  NAND2_X1 U2 ( .A1(n9), .A2(net223704), .ZN(net179236) );
  INV_X1 U3 ( .A(n8), .ZN(net223706) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(net240355) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n8) );
  CLKBUF_X1 U6 ( .A(n8), .Z(net241881) );
  CLKBUF_X1 U7 ( .A(B), .Z(n10) );
  NAND2_X1 U8 ( .A1(n10), .A2(A), .ZN(net223704) );
  XNOR2_X1 U9 ( .A(net240355), .B(net241881), .ZN(S) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  INV_X1 U2 ( .A(Ci), .ZN(n10) );
  NOR2_X1 U3 ( .A1(B), .A2(A), .ZN(n11) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n9) );
  OAI21_X1 U5 ( .B1(n11), .B2(n10), .A(n9), .ZN(Co) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n8), .S(S) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(n14), .Z(n9) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n13) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n14), .ZN(S) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n10) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n11) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n13) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n13), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n11), .B(n9), .ZN(S) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14, n15;

  CLKBUF_X1 U1 ( .A(n15), .Z(n9) );
  CLKBUF_X1 U2 ( .A(B), .Z(n10) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n11) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n15) );
  NAND2_X1 U5 ( .A1(n10), .A2(A), .ZN(n14) );
  INV_X1 U6 ( .A(n15), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n12), .A2(Ci), .ZN(n13) );
  NAND2_X1 U8 ( .A1(n13), .A2(n14), .ZN(Co) );
  XNOR2_X1 U9 ( .A(n11), .B(n9), .ZN(S) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net179251, n7, n8, n9, n10;
  assign Co = net179251;

  CLKBUF_X1 U1 ( .A(B), .Z(n7) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n10), .ZN(net179251) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NOR2_X1 U5 ( .A1(B), .A2(A), .ZN(n8) );
  FA_X1 U6 ( .A(n7), .B(A), .CI(Ci), .S(S) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(n9), .A2(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_15 UIV ( .A(S), .Y(SB) );
  ND2_45 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_44 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_43 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n10) );
  INV_X1 U4 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n9) );
  XNOR2_X1 U6 ( .A(n8), .B(n11), .ZN(S) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  BUF_X1 U1 ( .A(n10), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n11), .Z(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n10) );
  INV_X1 U5 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n9) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  OR2_X1 U2 ( .A1(n10), .A2(n13), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net179854, n8, n9, n10, n11, n12, n13;
  assign Co = net179854;

  XNOR2_X1 U1 ( .A(A), .B(Ci), .ZN(n12) );
  XNOR2_X1 U2 ( .A(n13), .B(n12), .ZN(S) );
  NAND2_X1 U3 ( .A1(A), .A2(Ci), .ZN(n11) );
  NOR2_X1 U4 ( .A1(A), .A2(Ci), .ZN(n10) );
  CLKBUF_X1 U5 ( .A(n9), .Z(n8) );
  OAI21_X1 U6 ( .B1(n9), .B2(n10), .A(n11), .ZN(net179854) );
  INV_X1 U7 ( .A(B), .ZN(n9) );
  INV_X1 U8 ( .A(n8), .ZN(n13) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(B), .Z(n9) );
  OAI21_X1 U2 ( .B1(n12), .B2(n11), .A(n10), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n11) );
  NOR2_X1 U4 ( .A1(B), .A2(A), .ZN(n12) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n10) );
  FA_X1 U6 ( .A(n9), .B(A), .CI(Ci), .S(S) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_53 UIV ( .A(S), .Y(SB) );
  ND2_159 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_158 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_157 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n8) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14, n15, n16;

  CLKBUF_X1 U1 ( .A(B), .Z(n10) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n11) );
  CLKBUF_X1 U3 ( .A(n16), .Z(n12) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n16) );
  NAND2_X1 U5 ( .A1(A), .A2(n10), .ZN(n15) );
  INV_X1 U6 ( .A(n12), .ZN(n13) );
  NAND2_X1 U7 ( .A1(n11), .A2(n13), .ZN(n14) );
  NAND2_X1 U8 ( .A1(n15), .A2(n14), .ZN(Co) );
  XNOR2_X1 U9 ( .A(Ci), .B(n16), .ZN(S) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  OAI21_X1 U1 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n10) );
  OR2_X1 U2 ( .A1(n11), .A2(n14), .ZN(n12) );
  INV_X1 U3 ( .A(n10), .ZN(n11) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n14) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n13) );
  NAND2_X1 U6 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n14), .ZN(S) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n13) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n9) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(B), .Z(n7) );
  INV_X1 U2 ( .A(Ci), .ZN(n9) );
  OAI21_X1 U3 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  NOR2_X1 U4 ( .A1(B), .A2(A), .ZN(n10) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n8) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n7), .S(S) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  INV_X1 U1 ( .A(n9), .ZN(n14) );
  INV_X1 U2 ( .A(A), .ZN(n10) );
  XNOR2_X1 U3 ( .A(n10), .B(B), .ZN(n9) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n13) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n9), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n11), .B(n14), .ZN(S) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net224803, n10, n11, n12, n13, n14;

  INV_X1 U1 ( .A(n11), .ZN(n13) );
  INV_X1 U2 ( .A(A), .ZN(n12) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U4 ( .A(B), .B(n12), .ZN(n11) );
  XNOR2_X1 U5 ( .A(n10), .B(n13), .ZN(S) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(net224803) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n11), .ZN(n14) );
  NAND2_X1 U8 ( .A1(n14), .A2(net224803), .ZN(Co) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  INV_X1 U1 ( .A(n10), .ZN(n13) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n9) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  INV_X1 U1 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n8) );
  OAI21_X1 U3 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  NOR2_X1 U4 ( .A1(B), .A2(A), .ZN(n10) );
  FA_X1 U5 ( .A(Ci), .B(A), .CI(B), .S(S) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n13) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U3 ( .A(n13), .ZN(n10) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U5 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_80 UIV ( .A(S), .Y(SB) );
  ND2_240 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_239 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_238 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n10) );
  INV_X1 U4 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n9) );
  XNOR2_X1 U6 ( .A(n8), .B(n11), .ZN(S) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(n9), .B(n13), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U5 ( .A(n13), .ZN(n10) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n12), .A2(n11), .ZN(Co) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net181057, net240110, net240360, net225339, net225338, n11, n12;
  assign Co = net181057;

  INV_X1 U1 ( .A(A), .ZN(n11) );
  XNOR2_X1 U2 ( .A(B), .B(n11), .ZN(n12) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n12), .ZN(net225339) );
  NAND2_X1 U4 ( .A1(net225339), .A2(net225338), .ZN(net181057) );
  INV_X1 U5 ( .A(n12), .ZN(net240360) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(net240110) );
  NAND2_X1 U7 ( .A1(B), .A2(A), .ZN(net225338) );
  XNOR2_X1 U8 ( .A(net240110), .B(net240360), .ZN(S) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net181060, n7, n8, n9, n10;
  assign Co = net181060;

  XNOR2_X1 U1 ( .A(A), .B(Ci), .ZN(n9) );
  XNOR2_X1 U2 ( .A(n10), .B(n9), .ZN(S) );
  NOR2_X1 U3 ( .A1(A), .A2(Ci), .ZN(n7) );
  AOI21_X1 U4 ( .B1(A), .B2(Ci), .A(B), .ZN(n8) );
  NOR2_X1 U5 ( .A1(n8), .A2(n7), .ZN(net181060) );
  CLKBUF_X1 U6 ( .A(B), .Z(n10) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net225353, net225355, net241877, n10, n11, n12, n13;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n10) );
  CLKBUF_X1 U2 ( .A(n10), .Z(net241877) );
  INV_X1 U3 ( .A(n10), .ZN(net225355) );
  CLKBUF_X1 U4 ( .A(B), .Z(n11) );
  NAND2_X1 U5 ( .A1(n11), .A2(A), .ZN(net225353) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n12) );
  NAND2_X1 U7 ( .A1(net225355), .A2(Ci), .ZN(n13) );
  NAND2_X1 U8 ( .A1(n13), .A2(net225353), .ZN(Co) );
  XNOR2_X1 U9 ( .A(n12), .B(net241877), .ZN(S) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  INV_X1 U2 ( .A(Ci), .ZN(n10) );
  NOR2_X1 U3 ( .A1(B), .A2(A), .ZN(n11) );
  OAI21_X1 U4 ( .B1(n11), .B2(n10), .A(n9), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n9) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n8), .S(S) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n11), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U6 ( .A(n9), .ZN(n13) );
  XNOR2_X1 U7 ( .A(n13), .B(n12), .ZN(S) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  CLKBUF_X1 U1 ( .A(n10), .Z(n8) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n10) );
  XOR2_X1 U3 ( .A(n8), .B(n11), .Z(S) );
  OAI21_X1 U4 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  INV_X1 U5 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n9) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n14) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n13) );
  INV_X1 U4 ( .A(n14), .ZN(n11) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n11), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n13), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n10), .B(n14), .ZN(S) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n10) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n14) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n13) );
  INV_X1 U4 ( .A(n14), .ZN(n11) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n11), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n10), .B(n14), .ZN(S) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XOR2_X1 U2 ( .A(n9), .B(n10), .Z(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U4 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n10) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  INV_X1 U3 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  INV_X1 U5 ( .A(n10), .ZN(n12) );
  XNOR2_X1 U6 ( .A(n12), .B(n11), .ZN(S) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(n8), .B(Ci), .ZN(S) );
  CLKBUF_X1 U2 ( .A(n10), .Z(n8) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n10) );
  OAI21_X1 U4 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  INV_X1 U5 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n9) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(n9), .Z(n7) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n9) );
  OAI21_X1 U3 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XOR2_X1 U4 ( .A(n7), .B(n10), .Z(S) );
  INV_X1 U5 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14, n15;

  CLKBUF_X1 U1 ( .A(n15), .Z(n10) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n11) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n15) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n14) );
  INV_X1 U5 ( .A(n15), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(Ci), .ZN(n13) );
  NAND2_X1 U7 ( .A1(n13), .A2(n14), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  INV_X1 U1 ( .A(Ci), .ZN(n9) );
  OAI21_X1 U2 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  NOR2_X1 U3 ( .A1(B), .A2(A), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  FA_X1 U5 ( .A(B), .B(A), .CI(Ci), .S(S) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net225936, net225938, n11, n12, n13;

  BUF_X1 U1 ( .A(n12), .Z(n11) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n12) );
  XNOR2_X1 U3 ( .A(Ci), .B(n11), .ZN(S) );
  INV_X1 U4 ( .A(n12), .ZN(net225938) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net225936) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net225938), .ZN(n13) );
  NAND2_X1 U7 ( .A1(n13), .A2(net225936), .ZN(Co) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(B), .Z(n7) );
  INV_X1 U2 ( .A(Ci), .ZN(n9) );
  OAI21_X1 U3 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n8) );
  NOR2_X1 U5 ( .A1(B), .A2(A), .ZN(n10) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n7), .S(S) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n11), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U6 ( .A(n9), .ZN(n13) );
  XNOR2_X1 U7 ( .A(n13), .B(n12), .ZN(S) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14;

  INV_X1 U1 ( .A(n10), .ZN(n14) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n10) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n13), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n11), .B(n14), .ZN(S) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  XNOR2_X1 U6 ( .A(n9), .B(n12), .ZN(S) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14, n15;

  CLKBUF_X1 U1 ( .A(n12), .Z(n10) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n11) );
  INV_X1 U3 ( .A(n10), .ZN(n15) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n12) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n14) );
  NAND2_X1 U6 ( .A1(n12), .A2(Ci), .ZN(n13) );
  NAND2_X1 U7 ( .A1(n13), .A2(n14), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n11), .B(n15), .ZN(S) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(B), .Z(n7) );
  INV_X1 U2 ( .A(Ci), .ZN(n9) );
  NOR2_X1 U3 ( .A1(B), .A2(A), .ZN(n10) );
  OAI21_X1 U4 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n8) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n7), .S(S) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(n11), .Z(n9) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n10) );
  XOR2_X1 U3 ( .A(n10), .B(n9), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n13) );
  NAND2_X1 U6 ( .A1(n11), .A2(Ci), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(Co) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(n12), .Z(n10) );
  OAI21_X1 U2 ( .B1(n12), .B2(n13), .A(n11), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n12) );
  INV_X1 U4 ( .A(Ci), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U6 ( .A(n10), .ZN(n14) );
  XNOR2_X1 U7 ( .A(n14), .B(n13), .ZN(S) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  BUF_X1 U1 ( .A(n11), .Z(n9) );
  OAI21_X1 U2 ( .B1(n11), .B2(n12), .A(n10), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n11) );
  INV_X1 U4 ( .A(Ci), .ZN(n12) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U6 ( .A(n9), .ZN(n13) );
  XNOR2_X1 U7 ( .A(n13), .B(n12), .ZN(S) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(n10), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n10) );
  OAI21_X1 U3 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n9) );
  INV_X1 U6 ( .A(n8), .ZN(n12) );
  XNOR2_X1 U7 ( .A(n12), .B(n11), .ZN(S) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  CLKBUF_X1 U1 ( .A(n10), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XOR2_X1 U3 ( .A(n8), .B(n11), .Z(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n10) );
  INV_X1 U5 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n9) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(B), .Z(n9) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(n9), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  OAI21_X1 U1 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n10) );
  INV_X1 U3 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  INV_X1 U5 ( .A(n10), .ZN(n12) );
  XNOR2_X1 U6 ( .A(n12), .B(n11), .ZN(S) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XOR2_X1 U1 ( .A(n8), .B(n9), .Z(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(n9), .B(n10), .Z(S) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U4 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14, n15;

  CLKBUF_X1 U1 ( .A(n10), .Z(n9) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n10) );
  INV_X1 U3 ( .A(n9), .ZN(n11) );
  CLKBUF_X1 U4 ( .A(B), .Z(n12) );
  CLKBUF_X1 U5 ( .A(Ci), .Z(n13) );
  NAND2_X1 U6 ( .A1(n12), .A2(A), .ZN(n15) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n10), .ZN(n14) );
  NAND2_X1 U8 ( .A1(n14), .A2(n15), .ZN(Co) );
  XNOR2_X1 U9 ( .A(n13), .B(n11), .ZN(S) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(B), .Z(n9) );
  INV_X1 U2 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n10) );
  NOR2_X1 U4 ( .A1(B), .A2(A), .ZN(n12) );
  OAI21_X1 U5 ( .B1(n12), .B2(n11), .A(n10), .ZN(Co) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n9), .S(S) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net182296, n8, n9, n10, n11, n12;
  assign Co = net182296;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n12) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n11), .ZN(n10) );
  NAND2_X1 U3 ( .A1(n10), .A2(n9), .ZN(net182296) );
  INV_X1 U4 ( .A(n8), .ZN(n11) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n8) );
  XNOR2_X1 U6 ( .A(n12), .B(n8), .ZN(S) );
  NAND2_X1 U7 ( .A1(A), .A2(B), .ZN(n9) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net182299, net241458, net241534, net226581, net226579, n10, n11, n12;
  assign Co = net182299;

  NAND2_X1 U1 ( .A1(net226581), .A2(Ci), .ZN(n11) );
  NAND2_X1 U2 ( .A1(n11), .A2(net226579), .ZN(net182299) );
  INV_X1 U3 ( .A(n10), .ZN(net226581) );
  CLKBUF_X1 U4 ( .A(Ci), .Z(net241534) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n10) );
  CLKBUF_X1 U6 ( .A(n10), .Z(net241458) );
  CLKBUF_X1 U7 ( .A(B), .Z(n12) );
  NAND2_X1 U8 ( .A1(A), .A2(n12), .ZN(net226579) );
  XNOR2_X1 U9 ( .A(net241534), .B(net241458), .ZN(S) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  OAI21_X1 U1 ( .B1(n10), .B2(n9), .A(n8), .ZN(Co) );
  CLKBUF_X1 U2 ( .A(B), .Z(n7) );
  INV_X1 U3 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n8) );
  NOR2_X1 U5 ( .A1(B), .A2(A), .ZN(n10) );
  FA_X1 U6 ( .A(Ci), .B(A), .CI(n7), .S(S) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9, n10;

  CLKBUF_X1 U1 ( .A(n9), .Z(n7) );
  XOR2_X1 U2 ( .A(n7), .B(n10), .Z(S) );
  OAI21_X1 U3 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U5 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n8) );
  OAI21_X1 U2 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n10) );
  INV_X1 U4 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n9) );
  XNOR2_X1 U6 ( .A(n8), .B(n11), .ZN(S) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n12) );
  INV_X1 U4 ( .A(n13), .ZN(n10) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(n9), .B(n10), .Z(S) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U4 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n8) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(n8), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n9) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(n8), .ZN(n12) );
  NAND2_X1 U5 ( .A1(n9), .A2(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n11), .A2(n12), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n10), .ZN(S) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  CLKBUF_X1 U1 ( .A(B), .Z(n8) );
  XOR2_X1 U2 ( .A(n10), .B(n11), .Z(S) );
  OAI21_X1 U3 ( .B1(n10), .B2(n11), .A(n9), .ZN(Co) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n10) );
  INV_X1 U5 ( .A(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(A), .A2(n8), .ZN(n9) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13, n14;

  CLKBUF_X1 U1 ( .A(n14), .Z(n10) );
  CLKBUF_X1 U2 ( .A(B), .Z(n9) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n14) );
  NAND2_X1 U4 ( .A1(A), .A2(n9), .ZN(n13) );
  INV_X1 U5 ( .A(n14), .ZN(n11) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n11), .ZN(n12) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n10), .ZN(S) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10;

  XOR2_X1 U1 ( .A(n9), .B(n10), .Z(S) );
  OAI21_X1 U2 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n9) );
  INV_X1 U4 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n8) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n9), .ZN(S) );
endmodule


module MUX21_212 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_212 UIV ( .A(S), .Y(SB) );
  ND2_636 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_635 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_634 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12, n13, n14;

  OAI21_X1 U1 ( .B1(n12), .B2(n13), .A(n11), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  INV_X1 U3 ( .A(Ci), .ZN(n13) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U5 ( .A(n12), .ZN(n14) );
  XNOR2_X1 U6 ( .A(n14), .B(n13), .ZN(S) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(Ci), .B(n12), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14;

  BUF_X1 U1 ( .A(n12), .Z(n10) );
  OAI21_X1 U2 ( .B1(n12), .B2(n13), .A(n11), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n12) );
  INV_X1 U4 ( .A(Ci), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U6 ( .A(n10), .ZN(n14) );
  XNOR2_X1 U7 ( .A(n14), .B(n13), .ZN(S) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(A), .Z(n8) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n9) );
  INV_X1 U3 ( .A(n10), .ZN(n13) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n10) );
  NAND2_X1 U5 ( .A1(n8), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n10), .ZN(n11) );
  NAND2_X1 U7 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n9), .B(n13), .ZN(S) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  INV_X1 U1 ( .A(n9), .ZN(n12) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n9) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n10), .A2(n11), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  INV_X1 U2 ( .A(Ci), .ZN(n8) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n7) );
  NOR2_X1 U4 ( .A1(A), .A2(B), .ZN(n9) );
  FA_X1 U5 ( .A(Ci), .B(B), .CI(A), .S(S) );
endmodule


module MUX21_220 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_220 UIV ( .A(S), .Y(SB) );
  ND2_660 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_659 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_658 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net227263, net227265, net241448, n9, n10;

  NAND2_X1 U1 ( .A1(Ci), .A2(net227265), .ZN(n10) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n9) );
  XNOR2_X1 U3 ( .A(net241448), .B(n9), .ZN(S) );
  INV_X1 U4 ( .A(n9), .ZN(net227265) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net227263) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(net241448) );
  NAND2_X1 U7 ( .A1(net227263), .A2(n10), .ZN(Co) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n10) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n13) );
  OAI21_X1 U4 ( .B1(n12), .B2(n13), .A(n11), .ZN(Co) );
  INV_X1 U5 ( .A(Ci), .ZN(n12) );
  XNOR2_X1 U6 ( .A(n13), .B(n10), .ZN(S) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n10, n11, n12, n13, n14, n15;

  CLKBUF_X1 U1 ( .A(A), .Z(n10) );
  INV_X1 U2 ( .A(B), .ZN(n11) );
  INV_X1 U3 ( .A(n11), .ZN(n12) );
  INV_X1 U4 ( .A(Ci), .ZN(n14) );
  OAI21_X1 U5 ( .B1(n15), .B2(n14), .A(n13), .ZN(Co) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n13) );
  NOR2_X1 U7 ( .A1(A), .A2(B), .ZN(n15) );
  FA_X1 U8 ( .A(Ci), .B(n10), .CI(n12), .S(S) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11, n12;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n8) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U4 ( .A(n12), .ZN(n9) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U6 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n8), .B(n12), .ZN(S) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n9) );
  XOR2_X1 U2 ( .A(n9), .B(Ci), .Z(S) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n10) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n12) );
  NAND2_X1 U5 ( .A1(n10), .A2(Ci), .ZN(n11) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11;

  INV_X1 U1 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n9) );
  NOR2_X1 U3 ( .A1(A), .A2(B), .ZN(n11) );
  OAI21_X1 U4 ( .B1(n11), .B2(n10), .A(n9), .ZN(Co) );
  FA_X1 U5 ( .A(Ci), .B(A), .CI(B), .S(S) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  INV_X1 U1 ( .A(Ci), .ZN(n8) );
  NOR2_X1 U2 ( .A1(A), .A2(B), .ZN(n9) );
  OAI21_X1 U3 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  FA_X1 U5 ( .A(Ci), .B(B), .CI(A), .S(S) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12, n13;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n9) );
  OR2_X1 U2 ( .A1(n10), .A2(n13), .ZN(n11) );
  INV_X1 U3 ( .A(n9), .ZN(n10) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n13) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n12) );
  NAND2_X1 U6 ( .A1(n12), .A2(n11), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n13), .ZN(S) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n9, n10, n11, n12;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n12) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n11) );
  INV_X1 U3 ( .A(n12), .ZN(n9) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n9), .ZN(n10) );
  NAND2_X1 U5 ( .A1(n11), .A2(n10), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n12), .ZN(S) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n11, n12, n13, n14, n15, n16, n17;

  BUF_X1 U1 ( .A(Ci), .Z(n12) );
  XNOR2_X1 U2 ( .A(n12), .B(n11), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n17) );
  INV_X1 U5 ( .A(A), .ZN(n14) );
  INV_X1 U6 ( .A(B), .ZN(n13) );
  NAND2_X1 U7 ( .A1(n14), .A2(n13), .ZN(n15) );
  NAND2_X1 U8 ( .A1(Ci), .A2(n15), .ZN(n16) );
  NAND2_X1 U9 ( .A1(n16), .A2(n17), .ZN(Co) );
endmodule


module FA_448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n9), .B2(n8), .A(n7), .ZN(Co) );
  INV_X1 U2 ( .A(Ci), .ZN(n8) );
  NOR2_X1 U3 ( .A1(A), .A2(B), .ZN(n9) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  FA_X1 U5 ( .A(A), .B(B), .CI(Ci), .S(S) );
endmodule


module FA_500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  OAI21_X1 U1 ( .B1(n9), .B2(n10), .A(n8), .ZN(Co) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n9) );
  INV_X1 U3 ( .A(Ci), .ZN(n10) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(n11) );
  XNOR2_X1 U6 ( .A(n11), .B(n10), .ZN(S) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  OAI21_X1 U1 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XOR2_X1 U2 ( .A(n8), .B(n9), .Z(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module FA_512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XOR2_X1 U1 ( .A(n8), .B(n9), .Z(S) );
  OAI21_X1 U2 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_4 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_3 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_2 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_1 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_16 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_15 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_14 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_13 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_20 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_19 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_18 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_17 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_6 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_24 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_23 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_22 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_21 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_9 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n2, n3, n4;
  assign n2 = S;

  MUX21_36 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n2), .Y(Y[0]) );
  MUX21_35 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n2), .Y(Y[1]) );
  MUX21_34 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_33 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n3), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n2), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n4), .Z(n3) );
endmodule


module RCA_gen_N4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_68 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_67 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_66 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_65 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_72 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_71 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_70 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_69 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_10 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_40 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_39 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_38 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_37 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_76 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_75 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_74 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_73 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_80 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_79 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_78 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_77 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_84 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_83 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_82 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_81 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_88 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_87 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_86 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_85 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_92 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_91 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_90 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_89 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_13 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_52 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_51 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_50 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_49 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_104 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_103 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_102 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_101 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_14 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_56 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_55 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_54 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_53 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_108 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_107 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_106 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_105 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_112 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_116 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_115 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_114 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_113 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_120 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_119 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_118 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_117 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_33 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_132 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_131 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_130 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_129 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_18 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_72 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_71 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_70 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_69 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_35 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_140 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_139 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_138 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_137 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_36 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_144 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_143 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_142 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_141 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_19 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_76 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_75 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_74 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_73 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_37 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_148 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_147 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_146 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_145 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_38 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_152 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_151 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_150 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_149 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_20 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_80 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_79 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_78 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_77 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_39 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_156 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_155 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_154 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_153 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_21 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_84 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_83 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_82 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_81 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_41 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_164 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_163 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_162 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_161 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_42 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_168 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_167 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_166 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_165 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_22 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_88 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_87 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_86 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_85 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_43 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_172 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_171 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_170 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_169 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_44 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_176 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_175 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_174 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_173 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_23 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_92 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_91 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_90 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_89 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_45 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_180 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_179 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_178 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_177 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_46 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_184 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_183 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_182 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_181 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_25 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;

  MUX21_100 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_99 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_98 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_97 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(S), .Z(n1) );
endmodule


module MUX21_GENERIC_N4_26 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2, n3;
  assign n1 = S;

  MUX21_104 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_103 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_102 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n3), .Y(Y[2]) );
  MUX21_101 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  BUF_X1 U1 ( .A(n1), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n1), .Z(n2) );
endmodule


module RCA_gen_N4_51 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_204 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_203 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_202 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_201 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_208 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_207 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_206 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_205 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_27 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;

  MUX21_108 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_107 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_106 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_105 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  BUF_X1 U1 ( .A(S), .Z(n1) );
endmodule


module RCA_gen_N4_53 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_212 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_211 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_210 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_209 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_216 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_215 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_214 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_213 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_28 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2, n3;
  assign n1 = S;

  MUX21_112 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_111 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_110 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_109 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n3), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n2) );
  CLKBUF_X1 U2 ( .A(n1), .Z(n3) );
endmodule


module RCA_gen_N4_55 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_220 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_219 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_218 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_217 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_224 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_223 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_222 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_221 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_29 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;
  assign n1 = S;

  MUX21_116 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_115 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_114 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_113 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
endmodule


module RCA_gen_N4_57 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_228 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_227 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_226 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_225 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_232 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_231 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_230 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_229 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_30 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;

  MUX21_120 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_119 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_118 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_117 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(S), .Z(n1) );
endmodule


module RCA_gen_N4_59 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_236 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_235 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_234 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_233 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_240 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_239 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_238 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_237 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_31 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_124 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_123 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_122 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_121 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_61 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_244 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_243 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_242 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_241 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_248 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_247 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_246 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_245 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_32 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_128 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_127 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_126 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_125 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_63 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_252 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_251 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_250 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_249 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_34 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_136 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_135 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_134 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_133 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  BUF_X1 U1 ( .A(n1), .Z(n2) );
endmodule


module MUX21_GENERIC_N4_35 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n2;
  assign n2 = S;

  MUX21_140 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n2), .Y(Y[0]) );
  MUX21_139 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n2), .Y(Y[1]) );
  MUX21_138 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_137 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
endmodule


module RCA_gen_N4_69 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_276 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_275 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_274 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_273 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_70 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_280 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_279 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_278 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_277 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_36 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;
  assign n1 = S;

  MUX21_144 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_143 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_142 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_141 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
endmodule


module RCA_gen_N4_71 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_284 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_283 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_282 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_281 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_72 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_288 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_287 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_286 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_285 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_37 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2, n3;
  assign n1 = S;

  MUX21_148 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_147 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_146 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n3), .Y(Y[2]) );
  MUX21_145 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n1), .Z(n2) );
endmodule


module RCA_gen_N4_73 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_292 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_291 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_290 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_289 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_74 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_296 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_295 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_294 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_293 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_38 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_152 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_151 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_150 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_149 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_75 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_300 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_299 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_298 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_297 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_76 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_304 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_303 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_302 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_301 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_39 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;
  assign n1 = S;

  MUX21_156 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_155 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_154 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_153 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
endmodule


module RCA_gen_N4_77 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_308 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_307 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_306 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_305 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_78 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_312 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_311 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_310 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_309 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_40 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_160 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_159 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_158 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_157 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_79 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_316 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_315 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_314 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_313 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_80 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_320 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_319 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_318 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_317 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_43 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;

  MUX21_172 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_171 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_170 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_169 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  BUF_X1 U1 ( .A(S), .Z(n1) );
  CLKBUF_X1 U2 ( .A(S), .Z(n2) );
endmodule


module RCA_gen_N4_85 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_340 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_339 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_338 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_337 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_86 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_344 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_343 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_342 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_341 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_44 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_176 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_175 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_174 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_173 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_87 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_348 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_347 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_346 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_345 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_88 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_352 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_351 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_350 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_349 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_45 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_180 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_179 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_178 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_177 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_89 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_356 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_355 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_354 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_353 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_90 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_360 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_359 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_358 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_357 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_46 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_184 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_183 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_182 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_181 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n2) );
endmodule


module RCA_gen_N4_91 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_364 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_363 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_362 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_361 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_92 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_368 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_367 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_366 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_365 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_47 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_188 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_187 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_186 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_185 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n2) );
endmodule


module RCA_gen_N4_93 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_372 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_371 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_370 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_369 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_94 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_376 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_375 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_374 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_373 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_48 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_192 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_191 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_190 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_189 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_95 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_380 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_379 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_378 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_377 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_96 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_384 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_383 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_382 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_381 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_51 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_204 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_203 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_202 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_201 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_102 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_408 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_407 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_406 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_405 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_52 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_208 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_207 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_206 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_205 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n2) );
endmodule


module MUX21_GENERIC_N4_53 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n2;
  assign n2 = S;

  MUX21_212 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n2), .Y(Y[0]) );
  MUX21_211 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n2), .Y(Y[1]) );
  MUX21_210 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_209 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
endmodule


module RCA_gen_N4_105 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_420 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_419 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_418 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_417 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_106 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_424 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_423 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_422 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_421 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_54 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1;
  assign n1 = S;

  MUX21_216 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_215 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_214 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_213 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
endmodule


module RCA_gen_N4_107 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_428 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_427 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_426 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_425 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_108 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_432 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_431 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_430 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_429 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_55 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;
  wire   n1, n2, n3;
  assign n1 = S;

  MUX21_220 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_219 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_218 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_217 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  INV_X1 U1 ( .A(n3), .ZN(n2) );
  INV_X1 U2 ( .A(n1), .ZN(n3) );
endmodule


module RCA_gen_N4_109 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_436 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_435 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_434 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_433 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_110 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_440 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_439 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_438 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_437 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_56 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_224 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_223 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_222 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_221 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_111 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_444 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_443 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_442 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_441 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_112 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_448 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_447 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_446 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_445 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_63 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_252 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_251 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_250 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_249 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_125 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_500 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_499 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_498 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_497 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_126 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_504 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_503 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_502 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_501 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_GENERIC_N4_0 ( A, B, S, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input S;


  MUX21_256 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_255 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_254 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_253 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
endmodule


module RCA_gen_N4_127 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_508 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_507 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_506 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_505 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_gen_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_512 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_511 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_510 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_509 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CSAdd_N4_1 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_2 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_1 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_1 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_2 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_4 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_3 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_2 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_3 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_6 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_5 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_3 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_4 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_8 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_7 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_4 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_5 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_10 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_9 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_5 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_6 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_12 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_11 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_6 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_7 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_14 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_13 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_7 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_4 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5;

  OR2_X2 U1 ( .A1(n5), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
endmodule


module genG_6 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genP_9 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  NAND2_X1 U1 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  AND2_X1 U4 ( .A1(P0), .A2(P1), .ZN(Pout) );
endmodule


module genG_8 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  INV_X1 U1 ( .A(G1), .ZN(n6) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
  NAND2_X2 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genP_20 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  OR2_X1 U2 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module CSAdd_N4_9 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_18 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_17 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_9 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_10 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_20 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_19 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_10 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_11 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_22 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_21 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_11 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_12 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_24 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_23 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_12 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_13 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_26 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_25 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_13 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_14 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_28 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_27 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_14 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_15 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_30 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_29 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_15 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_16 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_32 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_31 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_16 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_13 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genP_38 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  NAND2_X1 U2 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U3 ( .A(G1), .ZN(n8) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_43 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net180073, net238664, net224517, n6;
  assign Gout = net180073;
  assign Pout = net238664;

  NAND2_X1 U1 ( .A1(n6), .A2(net224517), .ZN(net180073) );
  INV_X1 U2 ( .A(G1), .ZN(net224517) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  AND2_X1 U4 ( .A1(P1), .A2(P0), .ZN(net238664) );
endmodule


module CSAdd_N4_17 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_34 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_33 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_17 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_18 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_36 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_35 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_18 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_19 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_38 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_37 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_19 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_20 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_40 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_39 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_20 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_21 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_42 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_41 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_21 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_22 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_44 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_43 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_22 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_23 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_46 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_45 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_23 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_24 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_48 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_47 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_24 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genP_64 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(G0), .A2(P1), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_65 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7;

  OR2_X2 U1 ( .A1(G1), .A2(n7), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_76 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module PGblock_71 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   net238538, n4;
  assign g = net238538;

  INV_X1 U1 ( .A(a), .ZN(n4) );
  XNOR2_X1 U2 ( .A(b), .B(n4), .ZN(p) );
  AND2_X1 U3 ( .A1(b), .A2(a), .ZN(net238538) );
endmodule


module PGblock_79 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n5;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n5) );
  XNOR2_X1 U3 ( .A(b), .B(n5), .ZN(p) );
endmodule


module PGblock_87 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4, n6;

  CLKBUF_X1 U1 ( .A(b), .Z(n4) );
  AND2_X1 U2 ( .A1(a), .A2(n4), .ZN(g) );
  INV_X1 U3 ( .A(a), .ZN(n6) );
  XNOR2_X1 U4 ( .A(b), .B(n6), .ZN(p) );
endmodule


module CSAdd_N4_25 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_50 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_49 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_25 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_26 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_52 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_51 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_26 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_27 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_54 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_53 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_27 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_28 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_56 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_55 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_28 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_29 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_58 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_57 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_29 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_30 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_60 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_59 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_30 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_31 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_62 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_61 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_31 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_32 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_64 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_63 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_32 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_31 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  INV_X1 U1 ( .A(n4), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
endmodule


module genP_90 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(n8), .A2(n7), .ZN(Gout) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genP_92 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  INV_X1 U1 ( .A(G1), .ZN(n8) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  NAND2_X1 U3 ( .A1(n8), .A2(n7), .ZN(Gout) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genG_35 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X2 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module genP_99 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module PGblock_103 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module CSAdd_N4_34 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_68 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_67 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_34 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_35 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_70 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_69 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_35 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_36 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_72 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_71 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_36 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_37 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_74 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_73 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_37 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_38 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_76 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_75 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_38 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_39 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_78 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_77 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_39 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_40 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_80 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_79 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_40 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_40 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net210570, n4, n5;
  assign Gout = net210570;

  OR2_X1 U1 ( .A1(G0), .A2(G1), .ZN(n4) );
  AND2_X2 U2 ( .A1(n4), .A2(n5), .ZN(net210570) );
  OR2_X1 U3 ( .A1(P1), .A2(G1), .ZN(n5) );
endmodule


module genG_42 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5;

  OR2_X2 U1 ( .A1(G1), .A2(n5), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
endmodule


module genP_112 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_120 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genG_45 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(P1), .A2(G0), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module PGblock_137 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_145 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3, n5;

  CLKBUF_X1 U1 ( .A(b), .Z(n3) );
  AND2_X1 U2 ( .A1(n3), .A2(a), .ZN(g) );
  INV_X1 U3 ( .A(a), .ZN(n5) );
  XNOR2_X1 U4 ( .A(b), .B(n5), .ZN(p) );
endmodule


module CSAdd_N4_42 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_84 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_83 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_42 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_43 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_86 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_85 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_43 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_44 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_88 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_87 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_44 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_45 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_90 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_89 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_45 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_46 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_92 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_91 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_46 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_47 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_94 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_93 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_47 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_48 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_96 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_95 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_48 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_49 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net213014, n5;
  assign Gout = net213014;

  OAI22_X1 U1 ( .A1(P1), .A2(G1), .B1(G0), .B2(G1), .ZN(n5) );
  INV_X1 U2 ( .A(n5), .ZN(net213014) );
endmodule


module genP_139 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6;

  OR2_X2 U1 ( .A1(G1), .A2(n6), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P0), .A2(P1), .ZN(Pout) );
  AND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
endmodule


module genG_52 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net182403, n4, n5;
  assign Gout = net182403;

  NAND2_X2 U1 ( .A1(n4), .A2(n5), .ZN(net182403) );
  NAND2_X1 U2 ( .A1(G0), .A2(P1), .ZN(n5) );
  INV_X1 U3 ( .A(G1), .ZN(n4) );
endmodule


module genP_145 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(G0), .A2(P1), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_157 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(Gout) );
endmodule


module PGblock_172 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_173 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_175 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_176 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module PGblock_184 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n5;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n5) );
  XNOR2_X1 U3 ( .A(b), .B(n5), .ZN(p) );
endmodule


module PGblock_185 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_186 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n4;

  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n4) );
  XNOR2_X1 U3 ( .A(b), .B(n4), .ZN(p) );
endmodule


module Gstart_6 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module CSAdd_N4_50 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_100 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_99 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_50 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_51 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_102 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_101 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_51 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_52 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_104 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_103 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_52 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_53 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_106 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_105 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_53 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_54 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_108 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_107 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_54 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_55 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_110 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_109 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_55 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_56 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_112 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_111 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_56 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_55 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(P1), .B2(G0), .A(G1), .ZN(n2) );
endmodule


module genG_58 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X2 U1 ( .A1(n5), .A2(n6), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n5) );
endmodule


module genP_163 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(P0), .ZN(Pout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module genG_59 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X2 U1 ( .A1(n4), .A2(G1), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genG_60 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net213703, n4;
  assign Gout = net213703;

  AOI21_X1 U1 ( .B1(G0), .B2(P1), .A(G1), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(net213703) );
endmodule


module genG_61 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net182991, net227340, n5;
  assign Gout = net182991;

  NAND2_X1 U1 ( .A1(G0), .A2(P1), .ZN(n5) );
  NAND2_X2 U2 ( .A1(n5), .A2(net227340), .ZN(net182991) );
  INV_X1 U3 ( .A(G1), .ZN(net227340) );
endmodule


module genP_168 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U2 ( .B1(G0), .B2(P1), .A(G1), .ZN(n2) );
  AND2_X1 U3 ( .A1(P1), .A2(P0), .ZN(Pout) );
endmodule


module genP_172 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_173 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genG_62 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   net183018, n4, n5;
  assign Gout = net183018;

  NAND2_X2 U1 ( .A1(n5), .A2(n4), .ZN(net183018) );
  INV_X1 U2 ( .A(G1), .ZN(n4) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n5) );
endmodule


module genP_176 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n2;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(n2), .ZN(Gout) );
  AOI21_X1 U3 ( .B1(G0), .B2(P1), .A(G1), .ZN(n2) );
endmodule


module genP_182 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_184 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(Gout) );
endmodule


module genP_185 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_187 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(Gout) );
endmodule


module genP_188 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P1), .A2(P0), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n6), .A2(n7), .ZN(Gout) );
endmodule


module genP_189 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   net183069, net233056, net227399, n6;
  assign Gout = net183069;
  assign Pout = net233056;

  NAND2_X1 U1 ( .A1(n6), .A2(net227399), .ZN(net183069) );
  INV_X1 U2 ( .A(G1), .ZN(net227399) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  AND2_X1 U4 ( .A1(P1), .A2(P0), .ZN(net233056) );
endmodule


module genG_63 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(G0), .A2(P1), .ZN(n5) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(Gout) );
endmodule


module PGblock_190 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PGblock_200 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_202 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_207 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3;

  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  INV_X1 U2 ( .A(a), .ZN(n3) );
  XNOR2_X1 U3 ( .A(b), .B(n3), .ZN(p) );
endmodule


module PGblock_210 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_211 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   n3, n4;

  CLKBUF_X1 U1 ( .A(a), .Z(n3) );
  CLKBUF_X1 U2 ( .A(b), .Z(n4) );
  AND2_X1 U3 ( .A1(n3), .A2(n4), .ZN(g) );
  XOR2_X1 U4 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_213 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(a), .B(b), .Z(p) );
endmodule


module PGblock_215 ( a, b, p, g );
  input a, b;
  output p, g;
  wire   net232863;

  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  CLKBUF_X1 U2 ( .A(a), .Z(net232863) );
  AND2_X1 U3 ( .A1(b), .A2(net232863), .ZN(g) );
endmodule


module PGblock_216 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module Gstart_7 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n7), .ZN(Gout) );
endmodule


module CSAdd_N4_63 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_126 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_125 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_63 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module CSAdd_N4_0 ( A, B, Ci, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;

  wire   [3:0] S1;
  wire   [3:0] S2;

  RCA_gen_N4_0 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S1) );
  RCA_gen_N4_127 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S2) );
  MUX21_GENERIC_N4_0 MUX ( .A(S1), .B(S2), .S(Ci), .Y(S) );
endmodule


module genG_69 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n4;

  OR2_X1 U1 ( .A1(G1), .A2(n4), .ZN(Gout) );
  AND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n4) );
endmodule


module genP_200 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  NAND2_X1 U2 ( .A1(n8), .A2(n7), .ZN(Gout) );
  INV_X1 U3 ( .A(G1), .ZN(n8) );
  NAND2_X1 U4 ( .A1(P1), .A2(G0), .ZN(n7) );
endmodule


module genG_71 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  NAND2_X1 U1 ( .A1(n6), .A2(n5), .ZN(Gout) );
  INV_X1 U2 ( .A(G1), .ZN(n6) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n5) );
endmodule


module genP_214 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n6, n7;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n7) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n6) );
  NAND2_X1 U4 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module genP_215 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genP_0 ( G1, P1, G0, P0, Pout, Gout );
  input G1, P1, G0, P0;
  output Pout, Gout;
  wire   n7, n8;

  AND2_X1 U1 ( .A1(P0), .A2(P1), .ZN(Pout) );
  INV_X1 U2 ( .A(G1), .ZN(n8) );
  NAND2_X1 U3 ( .A1(P1), .A2(G0), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n8), .A2(n7), .ZN(Gout) );
endmodule


module genG_0 ( G1, P1, G0, Gout );
  input G1, P1, G0;
  output Gout;
  wire   n5, n6;

  INV_X1 U1 ( .A(G1), .ZN(n6) );
  NAND2_X1 U2 ( .A1(P1), .A2(G0), .ZN(n5) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(Gout) );
endmodule


module PGblock_240 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module PGblock_247 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U1 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U2 ( .A1(a), .A2(b), .ZN(g) );
endmodule


module PGblock_0 ( a, b, p, g );
  input a, b;
  output p, g;


  AND2_X1 U1 ( .A1(a), .A2(b), .ZN(g) );
  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
endmodule


module Gstart_0 ( a, b, Cin, Gout );
  input a, b, Cin;
  output Gout;
  wire   n6, n7;

  NAND2_X1 U1 ( .A1(a), .A2(b), .ZN(n7) );
  OAI21_X1 U2 ( .B1(b), .B2(a), .A(Cin), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n7), .A2(n6), .ZN(Gout) );
endmodule


module SumGen_N32_1 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_8 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_7 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_6 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_5 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_4 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_3 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_2 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_1 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_1 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][24] , \GMat[2][20] , \GMat[2][16] , \GMat[2][12] ,
         \GMat[2][8] , \GMat[3][32] , \GMat[3][16] , \GMat[4][32] ,
         \GMat[4][28] , \PMat[0][32] , \PMat[0][31] , \PMat[0][30] ,
         \PMat[0][29] , \PMat[0][28] , \PMat[0][27] , \PMat[0][26] ,
         \PMat[0][25] , \PMat[0][24] , \PMat[0][23] , \PMat[0][22] ,
         \PMat[0][21] , \PMat[0][20] , \PMat[0][19] , \PMat[0][18] ,
         \PMat[0][17] , \PMat[0][16] , \PMat[0][15] , \PMat[0][14] ,
         \PMat[0][13] , \PMat[0][12] , \PMat[0][11] , \PMat[0][10] ,
         \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] , \PMat[0][5] ,
         \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][24] ,
         \PMat[2][20] , \PMat[2][16] , \PMat[2][12] , \PMat[2][8] ,
         \PMat[3][32] , \PMat[3][16] , \PMat[4][32] , \PMat[4][28] , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10;
  assign C[0] = Cin;
  assign C[4] = n3;

  Gstart_1 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_31 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_30 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_29 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_28 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_27 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_26 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_25 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_24 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_23 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_22 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_21 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_20 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_19 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_18 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_17 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_16 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_15 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_14 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_13 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_12 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_11 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_10 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_9 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_8 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_7 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_6 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_5 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_4 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_3 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_2 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_1 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_9 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_27 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_26 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_25 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_24 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_23 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), 
        .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_22 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), 
        .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_21 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), 
        .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_20 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), 
        .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_19 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(\GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(\GMat[1][20] ) );
  genP_18 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(\GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(\GMat[1][22] ) );
  genP_17 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(\GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(\GMat[1][24] ) );
  genP_16 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(\GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(\GMat[1][26] ) );
  genP_15 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(\GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(\GMat[1][28] ) );
  genP_14 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(\GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(\GMat[1][30] ) );
  genP_13 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(\GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(\GMat[1][32] ) );
  genG_8 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_12 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_11 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), 
        .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(\GMat[2][12] ) );
  genP_10 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), 
        .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_9 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), 
        .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(\GMat[2][20] ) );
  genP_8 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), 
        .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_7 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), 
        .P0(\PMat[1][26] ), .Pout(n1), .Gout(n2) );
  genP_6 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), 
        .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_7 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(C[2]) );
  genP_5 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(\GMat[2][12] ), 
        .P0(\PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_4 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(\GMat[2][20] ), 
        .P0(\PMat[2][20] ), .Pout(n4), .Gout(n5) );
  genP_3 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(n9), .P0(n10), 
        .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_6 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(\PMat[2][12] ), .G0(C[2]), .Gout(
        C[3]) );
  genG_5 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(C[2]), .Gout(n3) );
  genP_2 P2s_4_6 ( .G1(n2), .P1(n1), .G0(n5), .P0(n4), .Pout(\PMat[4][28] ), 
        .Gout(\GMat[4][28] ) );
  genP_1 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(n7), .P0(n8), 
        .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_4 G2s_5_4 ( .G1(\GMat[2][20] ), .P1(\PMat[2][20] ), .G0(n3), .Gout(C[5]) );
  genG_3 G2s_5_5 ( .G1(n5), .P1(n4), .G0(n6), .Gout(C[6]) );
  genG_2 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(n3), .Gout(C[7]) );
  genG_1 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n6), .Gout(C[8]) );
  BUF_X1 U1 ( .A(n3), .Z(n6) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n7) );
  CLKBUF_X1 U3 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U4 ( .A(n2), .Z(n9) );
  CLKBUF_X1 U5 ( .A(n1), .Z(n10) );
endmodule


module SumGen_N32_2 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_16 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_15 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_14 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_13 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_12 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_11 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_10 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_9 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_2 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][24] , \GMat[2][20] , \GMat[2][16] , \GMat[2][12] ,
         \GMat[2][8] , \GMat[3][32] , \GMat[3][16] , \GMat[4][32] ,
         \GMat[4][28] , \PMat[0][32] , \PMat[0][31] , \PMat[0][30] ,
         \PMat[0][29] , \PMat[0][28] , \PMat[0][27] , \PMat[0][26] ,
         \PMat[0][25] , \PMat[0][24] , \PMat[0][23] , \PMat[0][22] ,
         \PMat[0][21] , \PMat[0][20] , \PMat[0][19] , \PMat[0][18] ,
         \PMat[0][17] , \PMat[0][16] , \PMat[0][15] , \PMat[0][14] ,
         \PMat[0][13] , \PMat[0][12] , \PMat[0][11] , \PMat[0][10] ,
         \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] , \PMat[0][5] ,
         \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][24] ,
         \PMat[2][20] , \PMat[2][16] , \PMat[2][12] , \PMat[2][8] ,
         \PMat[3][32] , \PMat[3][16] , \PMat[4][32] , \PMat[4][28] , n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  assign C[0] = Cin;
  assign C[4] = n2;

  Gstart_2 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_62 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_61 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_60 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_59 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_58 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_57 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_56 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_55 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_54 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_53 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_52 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_51 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_50 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_49 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_48 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_47 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_46 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_45 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_44 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_43 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_42 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_41 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_40 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_39 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_38 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_37 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_36 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_35 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_34 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_33 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_32 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_18 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_54 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_53 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_52 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_51 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_50 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), 
        .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_49 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), 
        .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_48 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), 
        .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_47 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), 
        .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_46 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(\GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(\GMat[1][20] ) );
  genP_45 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(\GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(\GMat[1][22] ) );
  genP_44 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(\GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(\GMat[1][24] ) );
  genP_43 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(\GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(\GMat[1][26] ) );
  genP_42 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(\GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(\GMat[1][28] ) );
  genP_41 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(\GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(\GMat[1][30] ) );
  genP_40 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(\GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(\GMat[1][32] ) );
  genG_17 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_39 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_38 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), 
        .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(\GMat[2][12] ) );
  genP_37 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), 
        .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_36 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), 
        .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(\GMat[2][20] ) );
  genP_35 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), 
        .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_34 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), 
        .P0(\PMat[1][26] ), .Pout(n3), .Gout(n5) );
  genP_33 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), 
        .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_16 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(
        C[2]) );
  genP_32 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(\GMat[2][12] ), 
        .P0(\PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_31 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(\GMat[2][20] ), 
        .P0(\PMat[2][20] ), .Pout(n6), .Gout(n4) );
  genP_30 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(n12), .P0(n8), 
        .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_15 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(\PMat[2][12] ), .G0(C[2]), .Gout(
        C[3]) );
  genG_14 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(C[2]), .Gout(
        n2) );
  genP_29 P2s_4_6 ( .G1(n5), .P1(n3), .G0(n4), .P0(n11), .Pout(\PMat[4][28] ), 
        .Gout(\GMat[4][28] ) );
  genP_28 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(n10), .P0(n13), 
        .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_13 G2s_5_4 ( .G1(\GMat[2][20] ), .P1(\PMat[2][20] ), .G0(n2), .Gout(
        C[5]) );
  genG_12 G2s_5_5 ( .G1(n4), .P1(n6), .G0(n9), .Gout(C[6]) );
  genG_11 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(n7), .Gout(
        C[7]) );
  genG_10 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n7), .Gout(
        C[8]) );
  BUF_X1 U1 ( .A(n2), .Z(n9) );
  BUF_X1 U2 ( .A(n2), .Z(n7) );
  CLKBUF_X1 U3 ( .A(n3), .Z(n8) );
  CLKBUF_X1 U4 ( .A(n6), .Z(n11) );
  CLKBUF_X1 U5 ( .A(n4), .Z(n10) );
  CLKBUF_X1 U6 ( .A(n5), .Z(n12) );
  CLKBUF_X1 U7 ( .A(n11), .Z(n13) );
endmodule


module SumGen_N32_3 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_24 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_23 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_22 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_21 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_20 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_19 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_18 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_17 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_3 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][28] , \GMat[2][24] , \GMat[2][20] , \GMat[2][16] ,
         \GMat[2][12] , \GMat[2][8] , \GMat[3][32] , \GMat[3][16] ,
         \GMat[4][32] , \GMat[4][28] , \PMat[0][32] , \PMat[0][31] ,
         \PMat[0][30] , \PMat[0][29] , \PMat[0][28] , \PMat[0][27] ,
         \PMat[0][26] , \PMat[0][25] , \PMat[0][24] , \PMat[0][23] ,
         \PMat[0][22] , \PMat[0][21] , \PMat[0][20] , \PMat[0][19] ,
         \PMat[0][18] , \PMat[0][17] , \PMat[0][16] , \PMat[0][15] ,
         \PMat[0][14] , \PMat[0][13] , \PMat[0][12] , \PMat[0][11] ,
         \PMat[0][10] , \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] ,
         \PMat[0][5] , \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][24] ,
         \PMat[2][20] , \PMat[2][16] , \PMat[2][8] , \PMat[3][32] ,
         \PMat[3][16] , \PMat[4][32] , \PMat[4][28] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12;
  assign C[0] = Cin;
  assign C[4] = n4;

  Gstart_3 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_93 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_92 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_91 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_90 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_89 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_88 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_87 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_86 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_85 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_84 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_83 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_82 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_81 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_80 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_79 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_78 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_77 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_76 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_75 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_74 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_73 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_72 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_71 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_70 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_69 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_68 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_67 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_66 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_65 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_64 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_63 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_27 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_81 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_80 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_79 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_78 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_77 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), 
        .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_76 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), 
        .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_75 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), 
        .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_74 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), 
        .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_73 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(\GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(\GMat[1][20] ) );
  genP_72 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(\GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(\GMat[1][22] ) );
  genP_71 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(\GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(\GMat[1][24] ) );
  genP_70 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(\GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(\GMat[1][26] ) );
  genP_69 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(\GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(\GMat[1][28] ) );
  genP_68 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(\GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(\GMat[1][30] ) );
  genP_67 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(\GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(\GMat[1][32] ) );
  genG_26 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_66 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_65 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), 
        .P0(\PMat[1][10] ), .Pout(n1), .Gout(\GMat[2][12] ) );
  genP_64 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), 
        .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_63 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), 
        .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(\GMat[2][20] ) );
  genP_62 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), 
        .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_61 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), 
        .P0(\PMat[1][26] ), .Pout(n2), .Gout(\GMat[2][28] ) );
  genP_60 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), 
        .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_25 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(
        C[2]) );
  genP_59 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(\GMat[2][12] ), 
        .P0(n6), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_58 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(n10), .P0(
        \PMat[2][20] ), .Pout(n3), .Gout(n5) );
  genP_57 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(\GMat[2][28] ), 
        .P0(n11), .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_24 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(n1), .G0(C[2]), .Gout(C[3]) );
  genG_23 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(n7), .Gout(n4)
         );
  genP_56 P2s_4_6 ( .G1(\GMat[2][28] ), .P1(n2), .G0(n9), .P0(n12), .Pout(
        \PMat[4][28] ), .Gout(\GMat[4][28] ) );
  genP_55 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(n9), .P0(n12), 
        .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_22 G2s_5_4 ( .G1(\GMat[2][20] ), .P1(\PMat[2][20] ), .G0(n4), .Gout(
        C[5]) );
  genG_21 G2s_5_5 ( .G1(n5), .P1(n3), .G0(n8), .Gout(C[6]) );
  genG_20 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(n8), .Gout(
        C[7]) );
  genG_19 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n8), .Gout(
        C[8]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n6) );
  CLKBUF_X1 U2 ( .A(C[2]), .Z(n7) );
  CLKBUF_X1 U3 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U4 ( .A(n5), .Z(n9) );
  CLKBUF_X1 U5 ( .A(\GMat[2][20] ), .Z(n10) );
  CLKBUF_X1 U6 ( .A(n2), .Z(n11) );
  CLKBUF_X1 U7 ( .A(n3), .Z(n12) );
endmodule


module SumGen_N32_4 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_32 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_31 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_30 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_29 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_28 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_27 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_26 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_25 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_4 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][28] , \GMat[2][24] , \GMat[2][16] , \GMat[2][12] ,
         \GMat[2][8] , \GMat[3][32] , \GMat[3][16] , \GMat[4][32] ,
         \GMat[4][28] , \PMat[0][32] , \PMat[0][31] , \PMat[0][30] ,
         \PMat[0][29] , \PMat[0][28] , \PMat[0][27] , \PMat[0][26] ,
         \PMat[0][25] , \PMat[0][24] , \PMat[0][23] , \PMat[0][22] ,
         \PMat[0][21] , \PMat[0][20] , \PMat[0][19] , \PMat[0][18] ,
         \PMat[0][17] , \PMat[0][16] , \PMat[0][15] , \PMat[0][14] ,
         \PMat[0][13] , \PMat[0][12] , \PMat[0][11] , \PMat[0][10] ,
         \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] , \PMat[0][5] ,
         \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][24] ,
         \PMat[2][20] , \PMat[2][16] , \PMat[2][12] , \PMat[2][8] ,
         \PMat[3][32] , \PMat[3][16] , \PMat[4][32] , \PMat[4][28] , n1, n2,
         n3, n4, n5, n6, n7, n8;
  assign C[0] = Cin;
  assign C[4] = n3;

  Gstart_4 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_124 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_123 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_122 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_121 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_120 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_119 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_118 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_117 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_116 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_115 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_114 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_113 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_112 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_111 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_110 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_109 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_108 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_107 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_106 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_105 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_104 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_103 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_102 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_101 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_100 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_99 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_98 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_97 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_96 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_95 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_94 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_36 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_108 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_107 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_106 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_105 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_104 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_103 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_102 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_101 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_100 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(
        \GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(
        \GMat[1][20] ) );
  genP_99 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(\GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(\GMat[1][22] ) );
  genP_98 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(\GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(\GMat[1][24] ) );
  genP_97 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(\GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(\GMat[1][26] ) );
  genP_96 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(\GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(\GMat[1][28] ) );
  genP_95 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(\GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(\GMat[1][30] ) );
  genP_94 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(\GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(\GMat[1][32] ) );
  genG_35 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_93 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_92 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), 
        .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(\GMat[2][12] ) );
  genP_91 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), 
        .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_90 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), 
        .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(n4) );
  genP_89 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), 
        .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_88 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), 
        .P0(\PMat[1][26] ), .Pout(n1), .Gout(\GMat[2][28] ) );
  genP_87 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), 
        .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_34 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(
        C[2]) );
  genP_86 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(\GMat[2][12] ), 
        .P0(\PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_85 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(n4), .P0(
        \PMat[2][20] ), .Pout(n2), .Gout(n5) );
  genP_84 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(\GMat[2][28] ), 
        .P0(n1), .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_33 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(\PMat[2][12] ), .G0(C[2]), .Gout(
        C[3]) );
  genG_32 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(C[2]), .Gout(
        n3) );
  genP_83 P2s_4_6 ( .G1(\GMat[2][28] ), .P1(n1), .G0(n7), .P0(n8), .Pout(
        \PMat[4][28] ), .Gout(\GMat[4][28] ) );
  genP_82 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(n7), .P0(n8), 
        .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_31 G2s_5_4 ( .G1(n4), .P1(\PMat[2][20] ), .G0(n3), .Gout(C[5]) );
  genG_30 G2s_5_5 ( .G1(n5), .P1(n2), .G0(n3), .Gout(C[6]) );
  genG_29 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(n6), .Gout(
        C[7]) );
  genG_28 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n6), .Gout(
        C[8]) );
  CLKBUF_X1 U1 ( .A(n3), .Z(n6) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n7) );
  CLKBUF_X1 U3 ( .A(n2), .Z(n8) );
endmodule


module SumGen_N32_5 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_40 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_39 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_38 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_37 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_36 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_35 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_34 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_33 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_5 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][28] , \GMat[2][24] , \GMat[2][20] , \GMat[2][16] ,
         \GMat[2][8] , \GMat[3][32] , \GMat[3][16] , \GMat[4][32] ,
         \GMat[4][28] , \PMat[0][32] , \PMat[0][31] , \PMat[0][30] ,
         \PMat[0][29] , \PMat[0][28] , \PMat[0][27] , \PMat[0][26] ,
         \PMat[0][25] , \PMat[0][24] , \PMat[0][23] , \PMat[0][22] ,
         \PMat[0][21] , \PMat[0][20] , \PMat[0][19] , \PMat[0][18] ,
         \PMat[0][17] , \PMat[0][16] , \PMat[0][15] , \PMat[0][14] ,
         \PMat[0][13] , \PMat[0][12] , \PMat[0][11] , \PMat[0][10] ,
         \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] , \PMat[0][5] ,
         \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][28] ,
         \PMat[2][24] , \PMat[2][20] , \PMat[2][16] , \PMat[2][12] ,
         \PMat[2][8] , \PMat[3][32] , \PMat[3][16] , \PMat[4][32] ,
         \PMat[4][28] , n1, n2, n3, n4, n5, n7, n8, n9, n10;
  assign C[0] = Cin;
  assign C[4] = n5;

  Gstart_5 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_155 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_154 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_153 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_152 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_151 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_150 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_149 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_148 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_147 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_146 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_145 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_144 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_143 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_142 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_141 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_140 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_139 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_138 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_137 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_136 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_135 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_134 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_133 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_132 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_131 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_130 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_129 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_128 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_127 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_126 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_125 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_45 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_135 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_134 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_133 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_132 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_131 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_130 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_129 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_128 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_127 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(
        \GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(
        \GMat[1][20] ) );
  genP_126 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(
        \GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(
        \GMat[1][22] ) );
  genP_125 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(
        \GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(
        \GMat[1][24] ) );
  genP_124 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(
        \GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(
        \GMat[1][26] ) );
  genP_123 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(
        \GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(
        \GMat[1][28] ) );
  genP_122 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(
        \GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(
        \GMat[1][30] ) );
  genP_121 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(
        \GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(
        \GMat[1][32] ) );
  genG_44 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_120 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_119 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(n4) );
  genP_118 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_117 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(\GMat[2][20] ) );
  genP_116 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_115 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), .P0(\PMat[1][26] ), .Pout(\PMat[2][28] ), .Gout(\GMat[2][28] ) );
  genP_114 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_43 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(n1)
         );
  genP_113 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(n4), .P0(
        \PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_112 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(n8), .P0(
        \PMat[2][20] ), .Pout(n3), .Gout(n2) );
  genP_111 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(\GMat[2][28] ), .P0(\PMat[2][28] ), .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_42 G2s_4_2 ( .G1(n4), .P1(\PMat[2][12] ), .G0(n1), .Gout(C[3]) );
  genG_41 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(n7), .Gout(n5)
         );
  genP_110 P2s_4_6 ( .G1(\GMat[2][28] ), .P1(\PMat[2][28] ), .G0(n9), .P0(n3), 
        .Pout(\PMat[4][28] ), .Gout(\GMat[4][28] ) );
  genP_109 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(n9), .P0(n3), 
        .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_40 G2s_5_4 ( .G1(\GMat[2][20] ), .P1(\PMat[2][20] ), .G0(n5), .Gout(
        C[5]) );
  genG_39 G2s_5_5 ( .G1(n2), .P1(n3), .G0(n10), .Gout(C[6]) );
  genG_38 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(n10), .Gout(
        C[7]) );
  genG_37 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n10), .Gout(
        C[8]) );
  BUF_X2 U1 ( .A(n1), .Z(C[2]) );
  CLKBUF_X1 U2 ( .A(\GMat[2][20] ), .Z(n8) );
  CLKBUF_X1 U3 ( .A(C[2]), .Z(n7) );
  CLKBUF_X1 U4 ( .A(n2), .Z(n9) );
  CLKBUF_X1 U5 ( .A(n5), .Z(n10) );
endmodule


module SumGen_N32_6 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_48 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_47 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_46 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_45 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_44 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_43 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_42 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_41 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_6 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][28] , \GMat[2][24] , \GMat[2][20] , \GMat[2][16] ,
         \GMat[2][12] , \GMat[2][8] , \GMat[3][32] , \GMat[3][16] ,
         \GMat[4][32] , \GMat[4][28] , \PMat[0][32] , \PMat[0][31] ,
         \PMat[0][30] , \PMat[0][29] , \PMat[0][28] , \PMat[0][27] ,
         \PMat[0][26] , \PMat[0][25] , \PMat[0][24] , \PMat[0][23] ,
         \PMat[0][22] , \PMat[0][21] , \PMat[0][20] , \PMat[0][19] ,
         \PMat[0][18] , \PMat[0][17] , \PMat[0][16] , \PMat[0][15] ,
         \PMat[0][14] , \PMat[0][13] , \PMat[0][12] , \PMat[0][11] ,
         \PMat[0][10] , \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] ,
         \PMat[0][5] , \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][28] ,
         \PMat[2][24] , \PMat[2][20] , \PMat[2][16] , \PMat[2][12] ,
         \PMat[2][8] , \PMat[3][32] , \PMat[3][16] , \PMat[4][32] ,
         \PMat[4][28] , n1, n2, n3, n4, n5, n6, n7, n8;
  assign C[0] = Cin;
  assign C[2] = n2;
  assign C[4] = n4;

  Gstart_6 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_186 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_185 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_184 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_183 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_182 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_181 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_180 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_179 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_178 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_177 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_176 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_175 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_174 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_173 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_172 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_171 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_170 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_169 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_168 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_167 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_166 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_165 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_164 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_163 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_162 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_161 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_160 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_159 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_158 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_157 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_156 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_54 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_162 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_161 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_160 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_159 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_158 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_157 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_156 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_155 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_154 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(
        \GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(
        \GMat[1][20] ) );
  genP_153 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(
        \GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(
        \GMat[1][22] ) );
  genP_152 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(
        \GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(
        \GMat[1][24] ) );
  genP_151 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(
        \GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(
        \GMat[1][26] ) );
  genP_150 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(
        \GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(
        \GMat[1][28] ) );
  genP_149 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(
        \GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(
        \GMat[1][30] ) );
  genP_148 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(
        \GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(
        \GMat[1][32] ) );
  genG_53 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_147 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_146 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(\GMat[2][12] ) );
  genP_145 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_144 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(\GMat[2][20] ) );
  genP_143 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_142 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), .P0(\PMat[1][26] ), .Pout(\PMat[2][28] ), .Gout(\GMat[2][28] ) );
  genP_141 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_52 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(n2)
         );
  genP_140 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(n5), .P0(
        \PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_139 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(n6), .P0(
        \PMat[2][20] ), .Pout(n3), .Gout(n1) );
  genP_138 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(\GMat[2][28] ), .P0(\PMat[2][28] ), .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_51 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(\PMat[2][12] ), .G0(n2), .Gout(
        C[3]) );
  genG_50 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(n7), .Gout(n4)
         );
  genP_137 P2s_4_6 ( .G1(\GMat[2][28] ), .P1(\PMat[2][28] ), .G0(n1), .P0(n3), 
        .Pout(\PMat[4][28] ), .Gout(\GMat[4][28] ) );
  genP_136 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(n1), .P0(n3), 
        .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_49 G2s_5_4 ( .G1(\GMat[2][20] ), .P1(\PMat[2][20] ), .G0(n4), .Gout(
        C[5]) );
  genG_48 G2s_5_5 ( .G1(n1), .P1(n3), .G0(n4), .Gout(C[6]) );
  genG_47 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(n8), .Gout(
        C[7]) );
  genG_46 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n8), .Gout(
        C[8]) );
  CLKBUF_X1 U1 ( .A(\GMat[2][12] ), .Z(n5) );
  CLKBUF_X1 U2 ( .A(\GMat[2][20] ), .Z(n6) );
  CLKBUF_X1 U3 ( .A(n2), .Z(n7) );
  CLKBUF_X1 U4 ( .A(n4), .Z(n8) );
endmodule


module SumGen_N32_7 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_56 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_55 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_54 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_53 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_52 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_51 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_50 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_49 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_7 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][28] , \GMat[2][24] , \GMat[2][16] , \GMat[2][12] ,
         \GMat[2][8] , \GMat[3][32] , \GMat[3][24] , \GMat[3][16] ,
         \GMat[4][32] , \GMat[4][28] , \PMat[0][32] , \PMat[0][31] ,
         \PMat[0][30] , \PMat[0][29] , \PMat[0][28] , \PMat[0][27] ,
         \PMat[0][26] , \PMat[0][25] , \PMat[0][24] , \PMat[0][23] ,
         \PMat[0][22] , \PMat[0][21] , \PMat[0][20] , \PMat[0][19] ,
         \PMat[0][18] , \PMat[0][17] , \PMat[0][16] , \PMat[0][15] ,
         \PMat[0][14] , \PMat[0][13] , \PMat[0][12] , \PMat[0][11] ,
         \PMat[0][10] , \PMat[0][9] , \PMat[0][8] , \PMat[0][7] , \PMat[0][6] ,
         \PMat[0][5] , \PMat[0][4] , \PMat[0][3] , \PMat[0][2] , \PMat[1][32] ,
         \PMat[1][30] , \PMat[1][28] , \PMat[1][26] , \PMat[1][24] ,
         \PMat[1][22] , \PMat[1][20] , \PMat[1][18] , \PMat[1][16] ,
         \PMat[1][14] , \PMat[1][12] , \PMat[1][10] , \PMat[1][8] ,
         \PMat[1][6] , \PMat[1][4] , \PMat[2][32] , \PMat[2][28] ,
         \PMat[2][24] , \PMat[2][20] , \PMat[2][16] , \PMat[2][12] ,
         \PMat[2][8] , \PMat[3][32] , \PMat[3][24] , \PMat[3][16] ,
         \PMat[4][32] , \PMat[4][28] , n1, n2, n3, n4, n5;
  assign C[0] = Cin;
  assign C[2] = n1;

  Gstart_7 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_217 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_216 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_215 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_214 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_213 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_212 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_211 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_210 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_209 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_208 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_207 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_206 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_205 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_204 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_203 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_202 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_201 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_200 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_199 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_198 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_197 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_196 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_195 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_194 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_193 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_192 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_191 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_190 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_189 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_188 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_187 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_63 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_189 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_188 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_187 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_186 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_185 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_184 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_183 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_182 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_181 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(
        \GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(
        \GMat[1][20] ) );
  genP_180 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(
        \GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(
        \GMat[1][22] ) );
  genP_179 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(
        \GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(
        \GMat[1][24] ) );
  genP_178 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(
        \GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(
        \GMat[1][26] ) );
  genP_177 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(
        \GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(
        \GMat[1][28] ) );
  genP_176 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(
        \GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(
        \GMat[1][30] ) );
  genP_175 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(
        \GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(
        \GMat[1][32] ) );
  genG_62 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_174 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_173 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(\GMat[2][12] ) );
  genP_172 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_171 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(n2) );
  genP_170 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_169 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), .P0(\PMat[1][26] ), .Pout(\PMat[2][28] ), .Gout(\GMat[2][28] ) );
  genP_168 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_61 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(n1)
         );
  genP_167 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(n5), .P0(
        \PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_166 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(n2), .P0(
        \PMat[2][20] ), .Pout(\PMat[3][24] ), .Gout(\GMat[3][24] ) );
  genP_165 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(\GMat[2][28] ), .P0(\PMat[2][28] ), .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_60 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(\PMat[2][12] ), .G0(n1), .Gout(
        C[3]) );
  genG_59 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(n3), .Gout(
        C[4]) );
  genP_164 P2s_4_6 ( .G1(\GMat[2][28] ), .P1(\PMat[2][28] ), .G0(\GMat[3][24] ), .P0(\PMat[3][24] ), .Pout(\PMat[4][28] ), .Gout(\GMat[4][28] ) );
  genP_163 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(\GMat[3][24] ), .P0(\PMat[3][24] ), .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_58 G2s_5_4 ( .G1(n2), .P1(\PMat[2][20] ), .G0(C[4]), .Gout(C[5]) );
  genG_57 G2s_5_5 ( .G1(\GMat[3][24] ), .P1(\PMat[3][24] ), .G0(C[4]), .Gout(
        C[6]) );
  genG_56 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(C[4]), .Gout(
        C[7]) );
  genG_55 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(n4), .Gout(
        C[8]) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n3) );
  CLKBUF_X1 U2 ( .A(C[4]), .Z(n4) );
  CLKBUF_X1 U3 ( .A(\GMat[2][12] ), .Z(n5) );
endmodule


module SumGen_N32_0 ( A, B, C, S, Cout );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C;
  output [31:0] S;
  output Cout;

  assign Cout = C[8];

  CSAdd_N4_0 CSAs_0 ( .A(A[3:0]), .B(B[3:0]), .Ci(C[0]), .S(S[3:0]) );
  CSAdd_N4_63 CSAs_1 ( .A(A[7:4]), .B(B[7:4]), .Ci(C[1]), .S(S[7:4]) );
  CSAdd_N4_62 CSAs_2 ( .A(A[11:8]), .B(B[11:8]), .Ci(C[2]), .S(S[11:8]) );
  CSAdd_N4_61 CSAs_3 ( .A(A[15:12]), .B(B[15:12]), .Ci(C[3]), .S(S[15:12]) );
  CSAdd_N4_60 CSAs_4 ( .A(A[19:16]), .B(B[19:16]), .Ci(C[4]), .S(S[19:16]) );
  CSAdd_N4_59 CSAs_5 ( .A(A[23:20]), .B(B[23:20]), .Ci(C[5]), .S(S[23:20]) );
  CSAdd_N4_58 CSAs_6 ( .A(A[27:24]), .B(B[27:24]), .Ci(C[6]), .S(S[27:24]) );
  CSAdd_N4_57 CSAs_7 ( .A(A[31:28]), .B(B[31:28]), .Ci(C[7]), .S(S[31:28]) );
endmodule


module CarryGen_N32_0 ( A, B, Cin, C );
  input [32:1] A;
  input [32:1] B;
  output [8:0] C;
  input Cin;
  wire   Cin, \GMat[0][32] , \GMat[0][31] , \GMat[0][30] , \GMat[0][29] ,
         \GMat[0][28] , \GMat[0][27] , \GMat[0][26] , \GMat[0][25] ,
         \GMat[0][24] , \GMat[0][23] , \GMat[0][22] , \GMat[0][21] ,
         \GMat[0][20] , \GMat[0][19] , \GMat[0][18] , \GMat[0][17] ,
         \GMat[0][16] , \GMat[0][15] , \GMat[0][14] , \GMat[0][13] ,
         \GMat[0][12] , \GMat[0][11] , \GMat[0][10] , \GMat[0][9] ,
         \GMat[0][8] , \GMat[0][7] , \GMat[0][6] , \GMat[0][5] , \GMat[0][4] ,
         \GMat[0][3] , \GMat[0][2] , \GMat[0][1] , \GMat[1][32] ,
         \GMat[1][30] , \GMat[1][28] , \GMat[1][26] , \GMat[1][24] ,
         \GMat[1][22] , \GMat[1][20] , \GMat[1][18] , \GMat[1][16] ,
         \GMat[1][14] , \GMat[1][12] , \GMat[1][10] , \GMat[1][8] ,
         \GMat[1][6] , \GMat[1][4] , \GMat[1][2] , \GMat[2][32] ,
         \GMat[2][28] , \GMat[2][24] , \GMat[2][20] , \GMat[2][16] ,
         \GMat[2][12] , \GMat[2][8] , \GMat[3][32] , \GMat[3][24] ,
         \GMat[3][16] , \GMat[4][32] , \GMat[4][28] , \PMat[0][32] ,
         \PMat[0][31] , \PMat[0][30] , \PMat[0][29] , \PMat[0][28] ,
         \PMat[0][27] , \PMat[0][26] , \PMat[0][25] , \PMat[0][24] ,
         \PMat[0][23] , \PMat[0][22] , \PMat[0][21] , \PMat[0][20] ,
         \PMat[0][19] , \PMat[0][18] , \PMat[0][17] , \PMat[0][16] ,
         \PMat[0][15] , \PMat[0][14] , \PMat[0][13] , \PMat[0][12] ,
         \PMat[0][11] , \PMat[0][10] , \PMat[0][9] , \PMat[0][8] ,
         \PMat[0][7] , \PMat[0][6] , \PMat[0][5] , \PMat[0][4] , \PMat[0][3] ,
         \PMat[0][2] , \PMat[1][32] , \PMat[1][30] , \PMat[1][28] ,
         \PMat[1][26] , \PMat[1][24] , \PMat[1][22] , \PMat[1][20] ,
         \PMat[1][18] , \PMat[1][16] , \PMat[1][14] , \PMat[1][12] ,
         \PMat[1][10] , \PMat[1][8] , \PMat[1][6] , \PMat[1][4] ,
         \PMat[2][32] , \PMat[2][28] , \PMat[2][24] , \PMat[2][20] ,
         \PMat[2][16] , \PMat[2][12] , \PMat[2][8] , \PMat[3][32] ,
         \PMat[3][24] , \PMat[3][16] , \PMat[4][32] , \PMat[4][28] ;
  assign C[0] = Cin;

  Gstart_0 PG0_0_1 ( .a(A[1]), .b(B[1]), .Cin(Cin), .Gout(\GMat[0][1] ) );
  PGblock_0 PGs_0_2 ( .a(A[2]), .b(B[2]), .p(\PMat[0][2] ), .g(\GMat[0][2] )
         );
  PGblock_247 PGs_0_3 ( .a(A[3]), .b(B[3]), .p(\PMat[0][3] ), .g(\GMat[0][3] )
         );
  PGblock_246 PGs_0_4 ( .a(A[4]), .b(B[4]), .p(\PMat[0][4] ), .g(\GMat[0][4] )
         );
  PGblock_245 PGs_0_5 ( .a(A[5]), .b(B[5]), .p(\PMat[0][5] ), .g(\GMat[0][5] )
         );
  PGblock_244 PGs_0_6 ( .a(A[6]), .b(B[6]), .p(\PMat[0][6] ), .g(\GMat[0][6] )
         );
  PGblock_243 PGs_0_7 ( .a(A[7]), .b(B[7]), .p(\PMat[0][7] ), .g(\GMat[0][7] )
         );
  PGblock_242 PGs_0_8 ( .a(A[8]), .b(B[8]), .p(\PMat[0][8] ), .g(\GMat[0][8] )
         );
  PGblock_241 PGs_0_9 ( .a(A[9]), .b(B[9]), .p(\PMat[0][9] ), .g(\GMat[0][9] )
         );
  PGblock_240 PGs_0_10 ( .a(A[10]), .b(B[10]), .p(\PMat[0][10] ), .g(
        \GMat[0][10] ) );
  PGblock_239 PGs_0_11 ( .a(A[11]), .b(B[11]), .p(\PMat[0][11] ), .g(
        \GMat[0][11] ) );
  PGblock_238 PGs_0_12 ( .a(A[12]), .b(B[12]), .p(\PMat[0][12] ), .g(
        \GMat[0][12] ) );
  PGblock_237 PGs_0_13 ( .a(A[13]), .b(B[13]), .p(\PMat[0][13] ), .g(
        \GMat[0][13] ) );
  PGblock_236 PGs_0_14 ( .a(A[14]), .b(B[14]), .p(\PMat[0][14] ), .g(
        \GMat[0][14] ) );
  PGblock_235 PGs_0_15 ( .a(A[15]), .b(B[15]), .p(\PMat[0][15] ), .g(
        \GMat[0][15] ) );
  PGblock_234 PGs_0_16 ( .a(A[16]), .b(B[16]), .p(\PMat[0][16] ), .g(
        \GMat[0][16] ) );
  PGblock_233 PGs_0_17 ( .a(A[17]), .b(B[17]), .p(\PMat[0][17] ), .g(
        \GMat[0][17] ) );
  PGblock_232 PGs_0_18 ( .a(A[18]), .b(B[18]), .p(\PMat[0][18] ), .g(
        \GMat[0][18] ) );
  PGblock_231 PGs_0_19 ( .a(A[19]), .b(B[19]), .p(\PMat[0][19] ), .g(
        \GMat[0][19] ) );
  PGblock_230 PGs_0_20 ( .a(A[20]), .b(B[20]), .p(\PMat[0][20] ), .g(
        \GMat[0][20] ) );
  PGblock_229 PGs_0_21 ( .a(A[21]), .b(B[21]), .p(\PMat[0][21] ), .g(
        \GMat[0][21] ) );
  PGblock_228 PGs_0_22 ( .a(A[22]), .b(B[22]), .p(\PMat[0][22] ), .g(
        \GMat[0][22] ) );
  PGblock_227 PGs_0_23 ( .a(A[23]), .b(B[23]), .p(\PMat[0][23] ), .g(
        \GMat[0][23] ) );
  PGblock_226 PGs_0_24 ( .a(A[24]), .b(B[24]), .p(\PMat[0][24] ), .g(
        \GMat[0][24] ) );
  PGblock_225 PGs_0_25 ( .a(A[25]), .b(B[25]), .p(\PMat[0][25] ), .g(
        \GMat[0][25] ) );
  PGblock_224 PGs_0_26 ( .a(A[26]), .b(B[26]), .p(\PMat[0][26] ), .g(
        \GMat[0][26] ) );
  PGblock_223 PGs_0_27 ( .a(A[27]), .b(B[27]), .p(\PMat[0][27] ), .g(
        \GMat[0][27] ) );
  PGblock_222 PGs_0_28 ( .a(A[28]), .b(B[28]), .p(\PMat[0][28] ), .g(
        \GMat[0][28] ) );
  PGblock_221 PGs_0_29 ( .a(A[29]), .b(B[29]), .p(\PMat[0][29] ), .g(
        \GMat[0][29] ) );
  PGblock_220 PGs_0_30 ( .a(A[30]), .b(B[30]), .p(\PMat[0][30] ), .g(
        \GMat[0][30] ) );
  PGblock_219 PGs_0_31 ( .a(A[31]), .b(B[31]), .p(\PMat[0][31] ), .g(
        \GMat[0][31] ) );
  PGblock_218 PGs_0_32 ( .a(A[32]), .b(B[32]), .p(\PMat[0][32] ), .g(
        \GMat[0][32] ) );
  genG_0 G1s_1_1 ( .G1(\GMat[0][2] ), .P1(\PMat[0][2] ), .G0(\GMat[0][1] ), 
        .Gout(\GMat[1][2] ) );
  genP_0 P1s_1_2 ( .G1(\GMat[0][4] ), .P1(\PMat[0][4] ), .G0(\GMat[0][3] ), 
        .P0(\PMat[0][3] ), .Pout(\PMat[1][4] ), .Gout(\GMat[1][4] ) );
  genP_215 P1s_1_3 ( .G1(\GMat[0][6] ), .P1(\PMat[0][6] ), .G0(\GMat[0][5] ), 
        .P0(\PMat[0][5] ), .Pout(\PMat[1][6] ), .Gout(\GMat[1][6] ) );
  genP_214 P1s_1_4 ( .G1(\GMat[0][8] ), .P1(\PMat[0][8] ), .G0(\GMat[0][7] ), 
        .P0(\PMat[0][7] ), .Pout(\PMat[1][8] ), .Gout(\GMat[1][8] ) );
  genP_213 P1s_1_5 ( .G1(\GMat[0][10] ), .P1(\PMat[0][10] ), .G0(\GMat[0][9] ), 
        .P0(\PMat[0][9] ), .Pout(\PMat[1][10] ), .Gout(\GMat[1][10] ) );
  genP_212 P1s_1_6 ( .G1(\GMat[0][12] ), .P1(\PMat[0][12] ), .G0(\GMat[0][11] ), .P0(\PMat[0][11] ), .Pout(\PMat[1][12] ), .Gout(\GMat[1][12] ) );
  genP_211 P1s_1_7 ( .G1(\GMat[0][14] ), .P1(\PMat[0][14] ), .G0(\GMat[0][13] ), .P0(\PMat[0][13] ), .Pout(\PMat[1][14] ), .Gout(\GMat[1][14] ) );
  genP_210 P1s_1_8 ( .G1(\GMat[0][16] ), .P1(\PMat[0][16] ), .G0(\GMat[0][15] ), .P0(\PMat[0][15] ), .Pout(\PMat[1][16] ), .Gout(\GMat[1][16] ) );
  genP_209 P1s_1_9 ( .G1(\GMat[0][18] ), .P1(\PMat[0][18] ), .G0(\GMat[0][17] ), .P0(\PMat[0][17] ), .Pout(\PMat[1][18] ), .Gout(\GMat[1][18] ) );
  genP_208 P1s_1_10 ( .G1(\GMat[0][20] ), .P1(\PMat[0][20] ), .G0(
        \GMat[0][19] ), .P0(\PMat[0][19] ), .Pout(\PMat[1][20] ), .Gout(
        \GMat[1][20] ) );
  genP_207 P1s_1_11 ( .G1(\GMat[0][22] ), .P1(\PMat[0][22] ), .G0(
        \GMat[0][21] ), .P0(\PMat[0][21] ), .Pout(\PMat[1][22] ), .Gout(
        \GMat[1][22] ) );
  genP_206 P1s_1_12 ( .G1(\GMat[0][24] ), .P1(\PMat[0][24] ), .G0(
        \GMat[0][23] ), .P0(\PMat[0][23] ), .Pout(\PMat[1][24] ), .Gout(
        \GMat[1][24] ) );
  genP_205 P1s_1_13 ( .G1(\GMat[0][26] ), .P1(\PMat[0][26] ), .G0(
        \GMat[0][25] ), .P0(\PMat[0][25] ), .Pout(\PMat[1][26] ), .Gout(
        \GMat[1][26] ) );
  genP_204 P1s_1_14 ( .G1(\GMat[0][28] ), .P1(\PMat[0][28] ), .G0(
        \GMat[0][27] ), .P0(\PMat[0][27] ), .Pout(\PMat[1][28] ), .Gout(
        \GMat[1][28] ) );
  genP_203 P1s_1_15 ( .G1(\GMat[0][30] ), .P1(\PMat[0][30] ), .G0(
        \GMat[0][29] ), .P0(\PMat[0][29] ), .Pout(\PMat[1][30] ), .Gout(
        \GMat[1][30] ) );
  genP_202 P1s_1_16 ( .G1(\GMat[0][32] ), .P1(\PMat[0][32] ), .G0(
        \GMat[0][31] ), .P0(\PMat[0][31] ), .Pout(\PMat[1][32] ), .Gout(
        \GMat[1][32] ) );
  genG_71 G1s_2_1 ( .G1(\GMat[1][4] ), .P1(\PMat[1][4] ), .G0(\GMat[1][2] ), 
        .Gout(C[1]) );
  genP_201 P1s_2_2 ( .G1(\GMat[1][8] ), .P1(\PMat[1][8] ), .G0(\GMat[1][6] ), 
        .P0(\PMat[1][6] ), .Pout(\PMat[2][8] ), .Gout(\GMat[2][8] ) );
  genP_200 P1s_2_3 ( .G1(\GMat[1][12] ), .P1(\PMat[1][12] ), .G0(\GMat[1][10] ), .P0(\PMat[1][10] ), .Pout(\PMat[2][12] ), .Gout(\GMat[2][12] ) );
  genP_199 P1s_2_4 ( .G1(\GMat[1][16] ), .P1(\PMat[1][16] ), .G0(\GMat[1][14] ), .P0(\PMat[1][14] ), .Pout(\PMat[2][16] ), .Gout(\GMat[2][16] ) );
  genP_198 P1s_2_5 ( .G1(\GMat[1][20] ), .P1(\PMat[1][20] ), .G0(\GMat[1][18] ), .P0(\PMat[1][18] ), .Pout(\PMat[2][20] ), .Gout(\GMat[2][20] ) );
  genP_197 P1s_2_6 ( .G1(\GMat[1][24] ), .P1(\PMat[1][24] ), .G0(\GMat[1][22] ), .P0(\PMat[1][22] ), .Pout(\PMat[2][24] ), .Gout(\GMat[2][24] ) );
  genP_196 P1s_2_7 ( .G1(\GMat[1][28] ), .P1(\PMat[1][28] ), .G0(\GMat[1][26] ), .P0(\PMat[1][26] ), .Pout(\PMat[2][28] ), .Gout(\GMat[2][28] ) );
  genP_195 P1s_2_8 ( .G1(\GMat[1][32] ), .P1(\PMat[1][32] ), .G0(\GMat[1][30] ), .P0(\PMat[1][30] ), .Pout(\PMat[2][32] ), .Gout(\GMat[2][32] ) );
  genG_70 G2s_3_1 ( .G1(\GMat[2][8] ), .P1(\PMat[2][8] ), .G0(C[1]), .Gout(
        C[2]) );
  genP_194 P2s_3_3 ( .G1(\GMat[2][16] ), .P1(\PMat[2][16] ), .G0(\GMat[2][12] ), .P0(\PMat[2][12] ), .Pout(\PMat[3][16] ), .Gout(\GMat[3][16] ) );
  genP_193 P2s_3_5 ( .G1(\GMat[2][24] ), .P1(\PMat[2][24] ), .G0(\GMat[2][20] ), .P0(\PMat[2][20] ), .Pout(\PMat[3][24] ), .Gout(\GMat[3][24] ) );
  genP_192 P2s_3_7 ( .G1(\GMat[2][32] ), .P1(\PMat[2][32] ), .G0(\GMat[2][28] ), .P0(\PMat[2][28] ), .Pout(\PMat[3][32] ), .Gout(\GMat[3][32] ) );
  genG_69 G2s_4_2 ( .G1(\GMat[2][12] ), .P1(\PMat[2][12] ), .G0(C[2]), .Gout(
        C[3]) );
  genG_68 G2s_4_3 ( .G1(\GMat[3][16] ), .P1(\PMat[3][16] ), .G0(C[2]), .Gout(
        C[4]) );
  genP_191 P2s_4_6 ( .G1(\GMat[2][28] ), .P1(\PMat[2][28] ), .G0(\GMat[3][24] ), .P0(\PMat[3][24] ), .Pout(\PMat[4][28] ), .Gout(\GMat[4][28] ) );
  genP_190 P2s_4_7 ( .G1(\GMat[3][32] ), .P1(\PMat[3][32] ), .G0(\GMat[3][24] ), .P0(\PMat[3][24] ), .Pout(\PMat[4][32] ), .Gout(\GMat[4][32] ) );
  genG_67 G2s_5_4 ( .G1(\GMat[2][20] ), .P1(\PMat[2][20] ), .G0(C[4]), .Gout(
        C[5]) );
  genG_66 G2s_5_5 ( .G1(\GMat[3][24] ), .P1(\PMat[3][24] ), .G0(C[4]), .Gout(
        C[6]) );
  genG_65 G2s_5_6 ( .G1(\GMat[4][28] ), .P1(\PMat[4][28] ), .G0(C[4]), .Gout(
        C[7]) );
  genG_64 G2s_5_7 ( .G1(\GMat[4][32] ), .P1(\PMat[4][32] ), .G0(C[4]), .Gout(
        C[8]) );
endmodule


module ND2_1939 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2224 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X2 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2227 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_N32_1 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_288 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_287 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_286 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_285 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_284 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_283 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_282 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_281 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_280 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n5), .Y(Y[8]) );
  MUX21_279 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n5), .Y(Y[9]) );
  MUX21_278 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n5), .Y(Y[10]) );
  MUX21_277 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n5), .Y(Y[11]) );
  MUX21_276 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_275 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n4), .Y(Y[13]) );
  MUX21_274 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_273 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_272 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n4), .Y(Y[16]) );
  MUX21_271 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n4), .Y(Y[17]) );
  MUX21_270 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n4), .Y(Y[18]) );
  MUX21_269 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n6), .Y(Y[19]) );
  MUX21_268 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n6), .Y(Y[20]) );
  MUX21_267 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_266 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_265 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_264 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n5), .Y(Y[24]) );
  MUX21_263 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n5), .Y(Y[25]) );
  MUX21_262 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_261 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_260 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_259 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_258 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_257 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(n3), .Z(n6) );
  BUF_X1 U2 ( .A(n3), .Z(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n5) );
endmodule


module MUX21_GENERIC_N32_2 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n6, n7, n8, n9;
  assign n6 = S;

  MUX21_320 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n7), .Y(Y[0]) );
  MUX21_319 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n7), .Y(Y[1]) );
  MUX21_318 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n7), .Y(Y[2]) );
  MUX21_317 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n7), .Y(Y[3]) );
  MUX21_316 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n7), .Y(Y[4]) );
  MUX21_315 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n7), .Y(Y[5]) );
  MUX21_314 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n7), .Y(Y[6]) );
  MUX21_313 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n7), .Y(Y[7]) );
  MUX21_312 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n8), .Y(Y[8]) );
  MUX21_311 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n7), .Y(Y[9]) );
  MUX21_310 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n8), .Y(Y[10]) );
  MUX21_309 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n8), .Y(Y[11]) );
  MUX21_308 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n7), .Y(Y[12]) );
  MUX21_307 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n7), .Y(Y[13]) );
  MUX21_306 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n8), .Y(Y[14]) );
  MUX21_305 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n8), .Y(Y[15]) );
  MUX21_304 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n8), .Y(Y[16]) );
  MUX21_303 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n8), .Y(Y[17]) );
  MUX21_302 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n8), .Y(Y[18]) );
  MUX21_301 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n9), .Y(Y[19]) );
  MUX21_300 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n7), .Y(Y[20]) );
  MUX21_299 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n8), .Y(Y[21]) );
  MUX21_298 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n8), .Y(Y[22]) );
  MUX21_297 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n8), .Y(Y[23]) );
  MUX21_296 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n9), .Y(Y[24]) );
  MUX21_295 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n8), .Y(Y[25]) );
  MUX21_294 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n9), .Y(Y[26]) );
  MUX21_293 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n9), .Y(Y[27]) );
  MUX21_292 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n9), .Y(Y[28]) );
  MUX21_291 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n9), .Y(Y[29]) );
  MUX21_290 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n9), .Y(Y[30]) );
  MUX21_289 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n9), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(n6), .Z(n9) );
  BUF_X1 U2 ( .A(n6), .Z(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n7) );
endmodule


module MUX21_GENERIC_N32_5 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n5, n6, n7;
  assign n5 = S;

  MUX21_416 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n6), .Y(Y[0]) );
  MUX21_415 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n6), .Y(Y[1]) );
  MUX21_414 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n6), .Y(Y[2]) );
  MUX21_413 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n6), .Y(Y[3]) );
  MUX21_412 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n6), .Y(Y[4]) );
  MUX21_411 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n6), .Y(Y[5]) );
  MUX21_410 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n6), .Y(Y[6]) );
  MUX21_409 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n6), .Y(Y[7]) );
  MUX21_408 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n6), .Y(Y[8]) );
  MUX21_407 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n6), .Y(Y[9]) );
  MUX21_406 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n6), .Y(Y[10]) );
  MUX21_405 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n6), .Y(Y[11]) );
  MUX21_404 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n6), .Y(Y[12]) );
  MUX21_403 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n6), .Y(Y[13]) );
  MUX21_402 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n6), .Y(Y[14]) );
  MUX21_401 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n6), .Y(Y[15]) );
  MUX21_400 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n7), .Y(Y[16]) );
  MUX21_399 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n7), .Y(Y[17]) );
  MUX21_398 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n7), .Y(Y[18]) );
  MUX21_397 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n7), .Y(Y[19]) );
  MUX21_396 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n7), .Y(Y[20]) );
  MUX21_395 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n7), .Y(Y[21]) );
  MUX21_394 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n7), .Y(Y[22]) );
  MUX21_393 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n7), .Y(Y[23]) );
  MUX21_392 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n7), .Y(Y[24]) );
  MUX21_391 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n7), .Y(Y[25]) );
  MUX21_390 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n7), .Y(Y[26]) );
  MUX21_389 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n7), .Y(Y[27]) );
  MUX21_388 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n7), .Y(Y[28]) );
  MUX21_387 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n7), .Y(Y[29]) );
  MUX21_386 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n7), .Y(Y[30]) );
  MUX21_385 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n7), .Y(Y[31]) );
  BUF_X2 U1 ( .A(n5), .Z(n6) );
  BUF_X2 U2 ( .A(n5), .Z(n7) );
endmodule


module MUX21_GENERIC_N32_6 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n6, n7, n8, n9;
  assign n6 = S;

  MUX21_448 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n7), .Y(Y[0]) );
  MUX21_447 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n7), .Y(Y[1]) );
  MUX21_446 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n7), .Y(Y[2]) );
  MUX21_445 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n7), .Y(Y[3]) );
  MUX21_444 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n7), .Y(Y[4]) );
  MUX21_443 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n7), .Y(Y[5]) );
  MUX21_442 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n7), .Y(Y[6]) );
  MUX21_441 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n7), .Y(Y[7]) );
  MUX21_440 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n7), .Y(Y[8]) );
  MUX21_439 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n7), .Y(Y[9]) );
  MUX21_438 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n7), .Y(Y[10]) );
  MUX21_437 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n7), .Y(Y[11]) );
  MUX21_436 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n8), .Y(Y[12]) );
  MUX21_435 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n8), .Y(Y[13]) );
  MUX21_434 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n8), .Y(Y[14]) );
  MUX21_433 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n8), .Y(Y[15]) );
  MUX21_432 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n8), .Y(Y[16]) );
  MUX21_431 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n8), .Y(Y[17]) );
  MUX21_430 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n8), .Y(Y[18]) );
  MUX21_429 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n8), .Y(Y[19]) );
  MUX21_428 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n8), .Y(Y[20]) );
  MUX21_427 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n8), .Y(Y[21]) );
  MUX21_426 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n8), .Y(Y[22]) );
  MUX21_425 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n8), .Y(Y[23]) );
  MUX21_424 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n9), .Y(Y[24]) );
  MUX21_423 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n9), .Y(Y[25]) );
  MUX21_422 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n9), .Y(Y[26]) );
  MUX21_421 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n9), .Y(Y[27]) );
  MUX21_420 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n9), .Y(Y[28]) );
  MUX21_419 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n9), .Y(Y[29]) );
  MUX21_418 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n9), .Y(Y[30]) );
  MUX21_417 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n9), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n6), .Z(n7) );
  BUF_X1 U2 ( .A(n6), .Z(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n9) );
endmodule


module MUX21_GENERIC_N32_7 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n6, n7, n8;
  assign n6 = S;

  MUX21_480 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n7), .Y(Y[0]) );
  MUX21_479 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n8), .Y(Y[1]) );
  MUX21_478 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n8), .Y(Y[2]) );
  MUX21_477 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n8), .Y(Y[3]) );
  MUX21_476 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n8), .Y(Y[4]) );
  MUX21_475 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n8), .Y(Y[5]) );
  MUX21_474 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n8), .Y(Y[6]) );
  MUX21_473 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n8), .Y(Y[7]) );
  MUX21_472 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n8), .Y(Y[8]) );
  MUX21_471 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n8), .Y(Y[9]) );
  MUX21_470 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n8), .Y(Y[10]) );
  MUX21_469 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n8), .Y(Y[11]) );
  MUX21_468 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n8), .Y(Y[12]) );
  MUX21_467 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n8), .Y(Y[13]) );
  MUX21_466 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n8), .Y(Y[14]) );
  MUX21_465 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n7), .Y(Y[15]) );
  MUX21_464 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n8), .Y(Y[16]) );
  MUX21_463 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n7), .Y(Y[17]) );
  MUX21_462 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n7), .Y(Y[18]) );
  MUX21_461 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n7), .Y(Y[19]) );
  MUX21_460 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n7), .Y(Y[20]) );
  MUX21_459 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n7), .Y(Y[21]) );
  MUX21_458 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n7), .Y(Y[22]) );
  MUX21_457 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n7), .Y(Y[23]) );
  MUX21_456 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n7), .Y(Y[24]) );
  MUX21_455 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n7), .Y(Y[25]) );
  MUX21_454 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n7), .Y(Y[26]) );
  MUX21_453 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n7), .Y(Y[27]) );
  MUX21_452 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n7), .Y(Y[28]) );
  MUX21_451 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n7), .Y(Y[29]) );
  MUX21_450 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n7), .Y(Y[30]) );
  MUX21_449 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n8), .Y(Y[31]) );
  BUF_X2 U1 ( .A(n6), .Z(n7) );
  BUF_X2 U2 ( .A(n6), .Z(n8) );
endmodule


module Boothmul_N16_DW01_inc_6 ( A, SUM );
  input [32:0] A;
  output [32:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , n2;
  assign \carry[10]  = A[9];

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(\carry[11] ), .CO(\carry[12] ), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(n2), .CO(\carry[11] ), .S(SUM[10]) );
  XOR2_X1 U1_1_31 ( .A(A[31]), .B(\carry[31] ), .Z(SUM[31]) );
  INV_X1 U1 ( .A(SUM[9]), .ZN(n2) );
  INV_X1 U2 ( .A(\carry[10] ), .ZN(SUM[9]) );
endmodule


module Boothmul_N16_DW01_inc_5 ( A, SUM );
  input [32:0] A;
  output [32:0] SUM;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , n2;
  assign \carry[11]  = A[10];

  HA_X1 U1_1_30 ( .A(A[30]), .B(\carry[30] ), .CO(\carry[31] ), .S(SUM[30]) );
  HA_X1 U1_1_29 ( .A(A[29]), .B(\carry[29] ), .CO(\carry[30] ), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(\carry[28] ), .CO(\carry[29] ), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(\carry[27] ), .CO(\carry[28] ), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(\carry[26] ), .CO(\carry[27] ), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(\carry[25] ), .CO(\carry[26] ), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(\carry[24] ), .CO(\carry[25] ), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(\carry[23] ), .CO(\carry[24] ), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(\carry[22] ), .CO(\carry[23] ), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(\carry[21] ), .CO(\carry[22] ), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(\carry[20] ), .CO(\carry[21] ), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(\carry[19] ), .CO(\carry[20] ), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(\carry[18] ), .CO(\carry[19] ), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(\carry[17] ), .CO(\carry[18] ), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(\carry[16] ), .CO(\carry[17] ), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(\carry[15] ), .CO(\carry[16] ), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(\carry[14] ), .CO(\carry[15] ), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(\carry[13] ), .CO(\carry[14] ), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(\carry[12] ), .CO(\carry[13] ), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(n2), .CO(\carry[12] ), .S(SUM[11]) );
  XOR2_X1 U1_1_31 ( .A(A[31]), .B(\carry[31] ), .Z(SUM[31]) );
  INV_X1 U1 ( .A(SUM[10]), .ZN(n2) );
  INV_X1 U2 ( .A(\carry[11] ), .ZN(SUM[10]) );
endmodule


module p4adder_N32_1 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  wire   [8:0] C;
  assign n1 = B[11];
  assign n2 = B[15];
  assign n3 = B[19];
  assign n4 = B[28];
  assign n5 = B[23];
  assign n6 = B[27];
  assign n7 = B[31];
  assign n8 = B[30];

  CarryGen_N32_1 Cgen ( .A(A), .B({n12, n18, n19, n15, n6, B[26:24], n5, 
        B[22:20], n3, B[18:16], n2, B[14:12], n1, B[10:0]}), .Cin(Cin), .C(C)
         );
  SumGen_N32_1 Sgen ( .A(A), .B({n7, n8, B[29], n4, n17, n16, n20, B[24], n14, 
        B[22], n13, B[20], n3, B[18:16], n11, B[14:12], n9, B[10:8], n10, 
        B[6:0]}), .C(C), .S(S), .Cout(Cout) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n9) );
  BUF_X2 U2 ( .A(B[21]), .Z(n13) );
  CLKBUF_X1 U3 ( .A(B[7]), .Z(n10) );
  CLKBUF_X1 U4 ( .A(n2), .Z(n11) );
  BUF_X2 U5 ( .A(B[25]), .Z(n20) );
  CLKBUF_X1 U6 ( .A(n7), .Z(n12) );
  CLKBUF_X1 U7 ( .A(n5), .Z(n14) );
  CLKBUF_X1 U8 ( .A(n4), .Z(n15) );
  CLKBUF_X1 U9 ( .A(B[26]), .Z(n16) );
  CLKBUF_X1 U10 ( .A(n6), .Z(n17) );
  CLKBUF_X1 U11 ( .A(n8), .Z(n18) );
  CLKBUF_X1 U12 ( .A(B[29]), .Z(n19) );
endmodule


module mux51_generic_N32_1 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346;

  BUF_X4 U2 ( .A(n335), .Z(n233) );
  AND3_X1 U3 ( .A1(S[0]), .A2(S[1]), .A3(n242), .ZN(n225) );
  BUF_X4 U4 ( .A(n334), .Z(n231) );
  BUF_X1 U5 ( .A(n225), .Z(n230) );
  AND3_X1 U6 ( .A1(S[1]), .A2(n242), .A3(n244), .ZN(n226) );
  NAND2_X1 U7 ( .A1(n244), .A2(n241), .ZN(n343) );
  NAND3_X2 U8 ( .A1(n313), .A2(n312), .A3(n311), .ZN(Y[22]) );
  NAND3_X2 U9 ( .A1(n310), .A2(n309), .A3(n308), .ZN(Y[21]) );
  NAND3_X2 U10 ( .A1(n322), .A2(n321), .A3(n320), .ZN(Y[25]) );
  NAND3_X2 U11 ( .A1(n341), .A2(n340), .A3(n339), .ZN(Y[30]) );
  BUF_X2 U12 ( .A(n226), .Z(n236) );
  BUF_X2 U13 ( .A(n226), .Z(n235) );
  BUF_X2 U14 ( .A(n225), .Z(n228) );
  BUF_X2 U15 ( .A(n225), .Z(n229) );
  BUF_X2 U16 ( .A(n334), .Z(n232) );
  BUF_X2 U17 ( .A(n335), .Z(n234) );
  BUF_X2 U18 ( .A(n227), .Z(n238) );
  BUF_X2 U19 ( .A(n227), .Z(n237) );
  AND2_X1 U20 ( .A1(n244), .A2(n243), .ZN(n227) );
  AOI22_X1 U21 ( .A1(A[28]), .A2(n233), .B1(B[28]), .B2(n231), .ZN(n331) );
  NAND2_X1 U22 ( .A1(C[17]), .A2(n235), .ZN(n297) );
  AOI22_X1 U23 ( .A1(B[18]), .A2(n231), .B1(A[18]), .B2(n233), .ZN(n301) );
  AOI22_X1 U24 ( .A1(B[31]), .A2(n231), .B1(A[31]), .B2(n233), .ZN(n345) );
  NAND2_X1 U25 ( .A1(C[31]), .A2(n235), .ZN(n346) );
  AOI22_X1 U26 ( .A1(A[29]), .A2(n233), .B1(B[29]), .B2(n231), .ZN(n336) );
  AOI22_X1 U27 ( .A1(B[30]), .A2(n231), .B1(A[30]), .B2(n233), .ZN(n340) );
  NAND2_X1 U28 ( .A1(C[30]), .A2(n235), .ZN(n341) );
  AOI22_X1 U29 ( .A1(D[18]), .A2(n230), .B1(E[18]), .B2(n237), .ZN(n299) );
  NAND2_X1 U30 ( .A1(C[18]), .A2(n236), .ZN(n300) );
  NAND2_X1 U31 ( .A1(C[26]), .A2(n235), .ZN(n324) );
  NAND2_X1 U32 ( .A1(E[27]), .A2(n237), .ZN(n330) );
  AOI22_X1 U33 ( .A1(D[30]), .A2(n230), .B1(E[30]), .B2(n237), .ZN(n339) );
  NAND2_X1 U34 ( .A1(C[29]), .A2(n235), .ZN(n337) );
  AOI22_X1 U35 ( .A1(D[31]), .A2(n230), .B1(E[31]), .B2(n237), .ZN(n344) );
  AOI22_X1 U36 ( .A1(D[29]), .A2(n230), .B1(E[29]), .B2(n237), .ZN(n338) );
  NAND2_X1 U37 ( .A1(C[28]), .A2(n235), .ZN(n332) );
  AOI22_X1 U38 ( .A1(D[28]), .A2(n230), .B1(E[28]), .B2(n237), .ZN(n333) );
  INV_X1 U39 ( .A(B[27]), .ZN(n239) );
  INV_X1 U40 ( .A(S[2]), .ZN(n242) );
  INV_X1 U41 ( .A(S[1]), .ZN(n240) );
  NAND3_X1 U42 ( .A1(S[0]), .A2(n242), .A3(n240), .ZN(n342) );
  INV_X1 U43 ( .A(n342), .ZN(n334) );
  INV_X1 U44 ( .A(S[0]), .ZN(n244) );
  NOR2_X1 U45 ( .A1(S[2]), .A2(S[1]), .ZN(n241) );
  INV_X1 U46 ( .A(n343), .ZN(n335) );
  AOI22_X1 U47 ( .A1(B[0]), .A2(n232), .B1(A[0]), .B2(n234), .ZN(n247) );
  NAND2_X1 U48 ( .A1(C[0]), .A2(n236), .ZN(n246) );
  NOR2_X1 U49 ( .A1(n242), .A2(S[1]), .ZN(n243) );
  AOI22_X1 U50 ( .A1(D[0]), .A2(n228), .B1(E[0]), .B2(n238), .ZN(n245) );
  NAND3_X1 U51 ( .A1(n247), .A2(n246), .A3(n245), .ZN(Y[0]) );
  AOI22_X1 U52 ( .A1(B[1]), .A2(n232), .B1(A[1]), .B2(n234), .ZN(n250) );
  NAND2_X1 U53 ( .A1(C[1]), .A2(n235), .ZN(n249) );
  AOI22_X1 U54 ( .A1(D[1]), .A2(n228), .B1(E[1]), .B2(n237), .ZN(n248) );
  NAND3_X1 U55 ( .A1(n250), .A2(n249), .A3(n248), .ZN(Y[1]) );
  AOI22_X1 U56 ( .A1(B[2]), .A2(n232), .B1(A[2]), .B2(n234), .ZN(n253) );
  NAND2_X1 U57 ( .A1(C[2]), .A2(n236), .ZN(n252) );
  AOI22_X1 U58 ( .A1(D[2]), .A2(n228), .B1(E[2]), .B2(n238), .ZN(n251) );
  NAND3_X1 U59 ( .A1(n253), .A2(n252), .A3(n251), .ZN(Y[2]) );
  AOI22_X1 U60 ( .A1(B[3]), .A2(n232), .B1(A[3]), .B2(n234), .ZN(n256) );
  NAND2_X1 U61 ( .A1(C[3]), .A2(n236), .ZN(n255) );
  AOI22_X1 U62 ( .A1(D[3]), .A2(n228), .B1(E[3]), .B2(n238), .ZN(n254) );
  NAND3_X1 U63 ( .A1(n256), .A2(n255), .A3(n254), .ZN(Y[3]) );
  AOI22_X1 U64 ( .A1(B[4]), .A2(n232), .B1(A[4]), .B2(n234), .ZN(n259) );
  NAND2_X1 U65 ( .A1(C[4]), .A2(n236), .ZN(n258) );
  AOI22_X1 U66 ( .A1(D[4]), .A2(n228), .B1(E[4]), .B2(n238), .ZN(n257) );
  NAND3_X1 U67 ( .A1(n259), .A2(n258), .A3(n257), .ZN(Y[4]) );
  AOI22_X1 U68 ( .A1(B[5]), .A2(n232), .B1(A[5]), .B2(n234), .ZN(n262) );
  NAND2_X1 U69 ( .A1(C[5]), .A2(n236), .ZN(n261) );
  AOI22_X1 U70 ( .A1(D[5]), .A2(n228), .B1(E[5]), .B2(n238), .ZN(n260) );
  NAND3_X1 U71 ( .A1(n262), .A2(n261), .A3(n260), .ZN(Y[5]) );
  AOI22_X1 U72 ( .A1(B[6]), .A2(n232), .B1(A[6]), .B2(n234), .ZN(n265) );
  NAND2_X1 U73 ( .A1(C[6]), .A2(n236), .ZN(n264) );
  AOI22_X1 U74 ( .A1(D[6]), .A2(n228), .B1(E[6]), .B2(n238), .ZN(n263) );
  NAND3_X1 U75 ( .A1(n265), .A2(n264), .A3(n263), .ZN(Y[6]) );
  AOI22_X1 U76 ( .A1(B[7]), .A2(n232), .B1(A[7]), .B2(n234), .ZN(n268) );
  NAND2_X1 U77 ( .A1(C[7]), .A2(n236), .ZN(n267) );
  AOI22_X1 U78 ( .A1(D[7]), .A2(n228), .B1(E[7]), .B2(n238), .ZN(n266) );
  NAND3_X1 U79 ( .A1(n268), .A2(n267), .A3(n266), .ZN(Y[7]) );
  AOI22_X1 U80 ( .A1(B[8]), .A2(n232), .B1(A[8]), .B2(n234), .ZN(n271) );
  NAND2_X1 U81 ( .A1(C[8]), .A2(n236), .ZN(n270) );
  AOI22_X1 U82 ( .A1(D[8]), .A2(n228), .B1(E[8]), .B2(n238), .ZN(n269) );
  NAND3_X1 U83 ( .A1(n271), .A2(n270), .A3(n269), .ZN(Y[8]) );
  AOI22_X1 U84 ( .A1(B[9]), .A2(n231), .B1(A[9]), .B2(n233), .ZN(n274) );
  NAND2_X1 U85 ( .A1(C[9]), .A2(n236), .ZN(n273) );
  AOI22_X1 U86 ( .A1(D[9]), .A2(n228), .B1(E[9]), .B2(n238), .ZN(n272) );
  NAND3_X1 U87 ( .A1(n274), .A2(n273), .A3(n272), .ZN(Y[9]) );
  AOI22_X1 U88 ( .A1(B[10]), .A2(n231), .B1(A[10]), .B2(n233), .ZN(n277) );
  NAND2_X1 U89 ( .A1(C[10]), .A2(n236), .ZN(n276) );
  AOI22_X1 U90 ( .A1(D[10]), .A2(n228), .B1(E[10]), .B2(n238), .ZN(n275) );
  NAND3_X1 U91 ( .A1(n277), .A2(n276), .A3(n275), .ZN(Y[10]) );
  AOI22_X1 U92 ( .A1(B[11]), .A2(n231), .B1(A[11]), .B2(n233), .ZN(n280) );
  NAND2_X1 U93 ( .A1(C[11]), .A2(n236), .ZN(n279) );
  AOI22_X1 U94 ( .A1(D[11]), .A2(n228), .B1(E[11]), .B2(n238), .ZN(n278) );
  NAND3_X1 U95 ( .A1(n280), .A2(n279), .A3(n278), .ZN(Y[11]) );
  AOI22_X1 U96 ( .A1(B[12]), .A2(n231), .B1(A[12]), .B2(n233), .ZN(n283) );
  NAND2_X1 U97 ( .A1(C[12]), .A2(n236), .ZN(n282) );
  AOI22_X1 U98 ( .A1(D[12]), .A2(n229), .B1(E[12]), .B2(n238), .ZN(n281) );
  NAND3_X1 U99 ( .A1(n283), .A2(n282), .A3(n281), .ZN(Y[12]) );
  AOI22_X1 U100 ( .A1(B[13]), .A2(n231), .B1(A[13]), .B2(n233), .ZN(n286) );
  NAND2_X1 U101 ( .A1(C[13]), .A2(n236), .ZN(n285) );
  AOI22_X1 U102 ( .A1(D[13]), .A2(n229), .B1(E[13]), .B2(n238), .ZN(n284) );
  NAND3_X1 U103 ( .A1(n286), .A2(n285), .A3(n284), .ZN(Y[13]) );
  AOI22_X1 U104 ( .A1(B[14]), .A2(n231), .B1(A[14]), .B2(n233), .ZN(n289) );
  NAND2_X1 U105 ( .A1(C[14]), .A2(n236), .ZN(n288) );
  AOI22_X1 U106 ( .A1(D[14]), .A2(n229), .B1(E[14]), .B2(n238), .ZN(n287) );
  NAND3_X1 U107 ( .A1(n289), .A2(n288), .A3(n287), .ZN(Y[14]) );
  AOI22_X1 U108 ( .A1(B[15]), .A2(n231), .B1(A[15]), .B2(n233), .ZN(n292) );
  NAND2_X1 U109 ( .A1(C[15]), .A2(n236), .ZN(n291) );
  AOI22_X1 U110 ( .A1(D[15]), .A2(n229), .B1(E[15]), .B2(n238), .ZN(n290) );
  NAND3_X1 U111 ( .A1(n292), .A2(n291), .A3(n290), .ZN(Y[15]) );
  AOI22_X1 U112 ( .A1(B[16]), .A2(n231), .B1(A[16]), .B2(n233), .ZN(n295) );
  NAND2_X1 U113 ( .A1(C[16]), .A2(n235), .ZN(n294) );
  AOI22_X1 U114 ( .A1(D[16]), .A2(n229), .B1(E[16]), .B2(n238), .ZN(n293) );
  NAND3_X1 U115 ( .A1(n295), .A2(n294), .A3(n293), .ZN(Y[16]) );
  AOI22_X1 U116 ( .A1(B[17]), .A2(n231), .B1(A[17]), .B2(n233), .ZN(n298) );
  AOI22_X1 U117 ( .A1(D[17]), .A2(n229), .B1(E[17]), .B2(n237), .ZN(n296) );
  NAND3_X1 U118 ( .A1(n298), .A2(n297), .A3(n296), .ZN(Y[17]) );
  NAND3_X1 U119 ( .A1(n301), .A2(n300), .A3(n299), .ZN(Y[18]) );
  AOI22_X1 U120 ( .A1(B[19]), .A2(n231), .B1(A[19]), .B2(n233), .ZN(n304) );
  NAND2_X1 U121 ( .A1(C[19]), .A2(n235), .ZN(n303) );
  AOI22_X1 U122 ( .A1(D[19]), .A2(n229), .B1(E[19]), .B2(n237), .ZN(n302) );
  NAND3_X1 U123 ( .A1(n304), .A2(n303), .A3(n302), .ZN(Y[19]) );
  AOI22_X1 U124 ( .A1(B[20]), .A2(n231), .B1(A[20]), .B2(n233), .ZN(n307) );
  NAND2_X1 U125 ( .A1(C[20]), .A2(n235), .ZN(n306) );
  AOI22_X1 U126 ( .A1(D[20]), .A2(n229), .B1(E[20]), .B2(n237), .ZN(n305) );
  NAND3_X1 U127 ( .A1(n307), .A2(n306), .A3(n305), .ZN(Y[20]) );
  AOI22_X1 U128 ( .A1(B[21]), .A2(n231), .B1(A[21]), .B2(n233), .ZN(n310) );
  NAND2_X1 U129 ( .A1(C[21]), .A2(n235), .ZN(n309) );
  AOI22_X1 U130 ( .A1(D[21]), .A2(n229), .B1(E[21]), .B2(n237), .ZN(n308) );
  AOI22_X1 U131 ( .A1(B[22]), .A2(n231), .B1(A[22]), .B2(n233), .ZN(n313) );
  NAND2_X1 U132 ( .A1(C[22]), .A2(n235), .ZN(n312) );
  AOI22_X1 U133 ( .A1(D[22]), .A2(n229), .B1(E[22]), .B2(n237), .ZN(n311) );
  AOI22_X1 U134 ( .A1(B[23]), .A2(n231), .B1(A[23]), .B2(n233), .ZN(n316) );
  NAND2_X1 U135 ( .A1(C[23]), .A2(n235), .ZN(n315) );
  AOI22_X1 U136 ( .A1(D[23]), .A2(n229), .B1(E[23]), .B2(n237), .ZN(n314) );
  NAND3_X1 U137 ( .A1(n316), .A2(n315), .A3(n314), .ZN(Y[23]) );
  AOI22_X1 U138 ( .A1(B[24]), .A2(n231), .B1(A[24]), .B2(n233), .ZN(n319) );
  NAND2_X1 U139 ( .A1(C[24]), .A2(n235), .ZN(n318) );
  AOI22_X1 U140 ( .A1(D[24]), .A2(n229), .B1(E[24]), .B2(n237), .ZN(n317) );
  NAND3_X1 U141 ( .A1(n319), .A2(n318), .A3(n317), .ZN(Y[24]) );
  AOI22_X1 U142 ( .A1(B[25]), .A2(n231), .B1(A[25]), .B2(n233), .ZN(n322) );
  NAND2_X1 U143 ( .A1(C[25]), .A2(n235), .ZN(n321) );
  AOI22_X1 U144 ( .A1(D[25]), .A2(n230), .B1(E[25]), .B2(n237), .ZN(n320) );
  AOI22_X1 U145 ( .A1(B[26]), .A2(n231), .B1(A[26]), .B2(n233), .ZN(n325) );
  AOI22_X1 U146 ( .A1(D[26]), .A2(n230), .B1(E[26]), .B2(n237), .ZN(n323) );
  NAND3_X1 U147 ( .A1(n325), .A2(n324), .A3(n323), .ZN(Y[26]) );
  NAND2_X1 U148 ( .A1(D[27]), .A2(n230), .ZN(n329) );
  INV_X1 U149 ( .A(A[27]), .ZN(n326) );
  OAI22_X1 U150 ( .A1(n343), .A2(n326), .B1(n342), .B2(n239), .ZN(n327) );
  AOI21_X1 U151 ( .B1(C[27]), .B2(n235), .A(n327), .ZN(n328) );
  NAND3_X1 U152 ( .A1(n330), .A2(n329), .A3(n328), .ZN(Y[27]) );
  NAND3_X1 U153 ( .A1(n333), .A2(n332), .A3(n331), .ZN(Y[28]) );
  NAND3_X1 U154 ( .A1(n338), .A2(n337), .A3(n336), .ZN(Y[29]) );
  NAND3_X1 U155 ( .A1(n346), .A2(n345), .A3(n344), .ZN(Y[31]) );
endmodule


module p4adder_N32_2 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [8:0] C;
  assign n1 = B[7];
  assign n2 = B[11];
  assign n3 = B[29];
  assign n4 = B[28];
  assign n5 = B[26];
  assign n6 = B[23];
  assign n7 = B[27];

  CarryGen_N32_2 Cgen ( .A(A), .B({B[31:30], n14, n16, n7, n5, B[25:24], n6, 
        B[22:12], n2, B[10:8], n1, B[6:0]}), .Cin(Cin), .C(C) );
  SumGen_N32_2 Sgen ( .A(A), .B({B[31:30], n3, n4, n15, n9, B[25:24], n13, 
        B[22:20], n8, B[18:16], n12, B[14:12], n2, B[10:8], n11, B[6:4], n10, 
        B[2:0]}), .C(C), .S(S), .Cout(Cout) );
  CLKBUF_X1 U1 ( .A(B[19]), .Z(n8) );
  BUF_X2 U2 ( .A(n5), .Z(n9) );
  CLKBUF_X1 U3 ( .A(B[3]), .Z(n10) );
  CLKBUF_X1 U4 ( .A(n1), .Z(n11) );
  CLKBUF_X1 U5 ( .A(B[15]), .Z(n12) );
  CLKBUF_X1 U6 ( .A(n6), .Z(n13) );
  CLKBUF_X1 U7 ( .A(n3), .Z(n14) );
  CLKBUF_X1 U8 ( .A(n7), .Z(n15) );
  CLKBUF_X1 U9 ( .A(n4), .Z(n16) );
endmodule


module mux51_generic_N32_2 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351;

  INV_X2 U2 ( .A(n346), .ZN(n340) );
  INV_X2 U3 ( .A(n347), .ZN(n348) );
  INV_X2 U4 ( .A(n345), .ZN(n341) );
  AND3_X1 U5 ( .A1(S[1]), .A2(n242), .A3(n244), .ZN(n231) );
  NAND2_X1 U6 ( .A1(n244), .A2(n241), .ZN(n346) );
  NAND3_X4 U7 ( .A1(n283), .A2(n282), .A3(n281), .ZN(Y[12]) );
  NAND3_X2 U8 ( .A1(n335), .A2(n334), .A3(n333), .ZN(Y[28]) );
  BUF_X4 U9 ( .A(n231), .Z(n236) );
  BUF_X2 U10 ( .A(n231), .Z(n235) );
  BUF_X2 U11 ( .A(n329), .Z(n234) );
  BUF_X2 U12 ( .A(n232), .Z(n238) );
  BUF_X2 U13 ( .A(n232), .Z(n237) );
  INV_X1 U14 ( .A(n345), .ZN(n336) );
  AND2_X1 U15 ( .A1(n244), .A2(n243), .ZN(n232) );
  NAND2_X1 U16 ( .A1(C[15]), .A2(n235), .ZN(n291) );
  AOI22_X1 U17 ( .A1(B[29]), .A2(n336), .B1(A[29]), .B2(n340), .ZN(n338) );
  NAND2_X1 U18 ( .A1(C[29]), .A2(n235), .ZN(n339) );
  AOI22_X1 U19 ( .A1(D[29]), .A2(n348), .B1(E[29]), .B2(n237), .ZN(n337) );
  AOI22_X1 U20 ( .A1(B[30]), .A2(n341), .B1(A[30]), .B2(n340), .ZN(n343) );
  NAND2_X1 U21 ( .A1(C[30]), .A2(n235), .ZN(n344) );
  AOI22_X1 U22 ( .A1(D[30]), .A2(n348), .B1(E[30]), .B2(n237), .ZN(n342) );
  AOI22_X1 U23 ( .A1(B[31]), .A2(n336), .B1(A[31]), .B2(n340), .ZN(n350) );
  NAND2_X1 U24 ( .A1(C[31]), .A2(n235), .ZN(n351) );
  AOI22_X1 U25 ( .A1(D[31]), .A2(n348), .B1(E[31]), .B2(n237), .ZN(n349) );
  AOI22_X1 U26 ( .A1(A[26]), .A2(n340), .B1(B[26]), .B2(n341), .ZN(n326) );
  AOI22_X1 U27 ( .A1(B[28]), .A2(n336), .B1(A[28]), .B2(n340), .ZN(n334) );
  NAND2_X1 U28 ( .A1(C[28]), .A2(n235), .ZN(n335) );
  AOI22_X1 U29 ( .A1(A[27]), .A2(n340), .B1(B[27]), .B2(n341), .ZN(n330) );
  AOI22_X1 U30 ( .A1(B[16]), .A2(n341), .B1(A[16]), .B2(n340), .ZN(n295) );
  AOI22_X1 U31 ( .A1(D[16]), .A2(n348), .B1(E[16]), .B2(n237), .ZN(n293) );
  NAND2_X1 U32 ( .A1(C[16]), .A2(n235), .ZN(n294) );
  NAND2_X1 U33 ( .A1(C[24]), .A2(n235), .ZN(n318) );
  NAND2_X1 U34 ( .A1(E[25]), .A2(n237), .ZN(n325) );
  AOI22_X1 U35 ( .A1(D[28]), .A2(n348), .B1(E[28]), .B2(n237), .ZN(n333) );
  NAND2_X1 U36 ( .A1(C[27]), .A2(n235), .ZN(n331) );
  AOI22_X1 U37 ( .A1(D[27]), .A2(n348), .B1(E[27]), .B2(n237), .ZN(n332) );
  NAND2_X1 U38 ( .A1(C[26]), .A2(n235), .ZN(n327) );
  AOI22_X1 U39 ( .A1(D[26]), .A2(n348), .B1(E[26]), .B2(n237), .ZN(n328) );
  CLKBUF_X3 U40 ( .A(n320), .Z(n233) );
  INV_X1 U41 ( .A(B[25]), .ZN(n239) );
  INV_X1 U42 ( .A(S[2]), .ZN(n242) );
  INV_X1 U43 ( .A(S[1]), .ZN(n240) );
  NAND3_X1 U44 ( .A1(S[0]), .A2(n242), .A3(n240), .ZN(n345) );
  INV_X1 U45 ( .A(S[0]), .ZN(n244) );
  NOR2_X1 U46 ( .A1(S[2]), .A2(S[1]), .ZN(n241) );
  INV_X1 U47 ( .A(n346), .ZN(n329) );
  AOI22_X1 U48 ( .A1(B[0]), .A2(n341), .B1(A[0]), .B2(n234), .ZN(n247) );
  NAND2_X1 U49 ( .A1(C[0]), .A2(n236), .ZN(n246) );
  NAND3_X1 U50 ( .A1(S[0]), .A2(S[1]), .A3(n242), .ZN(n347) );
  INV_X1 U51 ( .A(n347), .ZN(n320) );
  NOR2_X1 U52 ( .A1(n242), .A2(S[1]), .ZN(n243) );
  AOI22_X1 U53 ( .A1(D[0]), .A2(n233), .B1(E[0]), .B2(n238), .ZN(n245) );
  NAND3_X1 U54 ( .A1(n247), .A2(n246), .A3(n245), .ZN(Y[0]) );
  AOI22_X1 U55 ( .A1(B[1]), .A2(n336), .B1(A[1]), .B2(n234), .ZN(n250) );
  NAND2_X1 U56 ( .A1(C[1]), .A2(n235), .ZN(n249) );
  AOI22_X1 U57 ( .A1(D[1]), .A2(n233), .B1(E[1]), .B2(n237), .ZN(n248) );
  NAND3_X1 U58 ( .A1(n250), .A2(n249), .A3(n248), .ZN(Y[1]) );
  AOI22_X1 U59 ( .A1(B[2]), .A2(n341), .B1(A[2]), .B2(n234), .ZN(n253) );
  NAND2_X1 U60 ( .A1(C[2]), .A2(n236), .ZN(n252) );
  AOI22_X1 U61 ( .A1(D[2]), .A2(n233), .B1(E[2]), .B2(n238), .ZN(n251) );
  NAND3_X1 U62 ( .A1(n253), .A2(n252), .A3(n251), .ZN(Y[2]) );
  AOI22_X1 U63 ( .A1(B[3]), .A2(n336), .B1(A[3]), .B2(n234), .ZN(n256) );
  NAND2_X1 U64 ( .A1(C[3]), .A2(n236), .ZN(n255) );
  AOI22_X1 U65 ( .A1(D[3]), .A2(n233), .B1(E[3]), .B2(n238), .ZN(n254) );
  NAND3_X1 U66 ( .A1(n256), .A2(n255), .A3(n254), .ZN(Y[3]) );
  AOI22_X1 U67 ( .A1(B[4]), .A2(n341), .B1(A[4]), .B2(n234), .ZN(n259) );
  NAND2_X1 U68 ( .A1(C[4]), .A2(n236), .ZN(n258) );
  AOI22_X1 U69 ( .A1(D[4]), .A2(n233), .B1(E[4]), .B2(n238), .ZN(n257) );
  NAND3_X1 U70 ( .A1(n259), .A2(n258), .A3(n257), .ZN(Y[4]) );
  AOI22_X1 U71 ( .A1(B[5]), .A2(n336), .B1(A[5]), .B2(n234), .ZN(n262) );
  NAND2_X1 U72 ( .A1(C[5]), .A2(n236), .ZN(n261) );
  AOI22_X1 U73 ( .A1(D[5]), .A2(n233), .B1(E[5]), .B2(n238), .ZN(n260) );
  NAND3_X1 U74 ( .A1(n262), .A2(n261), .A3(n260), .ZN(Y[5]) );
  AOI22_X1 U75 ( .A1(B[6]), .A2(n341), .B1(A[6]), .B2(n234), .ZN(n265) );
  NAND2_X1 U76 ( .A1(C[6]), .A2(n236), .ZN(n264) );
  AOI22_X1 U77 ( .A1(D[6]), .A2(n233), .B1(E[6]), .B2(n238), .ZN(n263) );
  NAND3_X1 U78 ( .A1(n265), .A2(n264), .A3(n263), .ZN(Y[6]) );
  AOI22_X1 U79 ( .A1(B[7]), .A2(n341), .B1(A[7]), .B2(n340), .ZN(n268) );
  NAND2_X1 U80 ( .A1(C[7]), .A2(n236), .ZN(n267) );
  AOI22_X1 U81 ( .A1(D[7]), .A2(n233), .B1(E[7]), .B2(n238), .ZN(n266) );
  NAND3_X1 U82 ( .A1(n268), .A2(n267), .A3(n266), .ZN(Y[7]) );
  AOI22_X1 U83 ( .A1(B[8]), .A2(n341), .B1(A[8]), .B2(n340), .ZN(n271) );
  NAND2_X1 U84 ( .A1(C[8]), .A2(n236), .ZN(n270) );
  AOI22_X1 U85 ( .A1(D[8]), .A2(n233), .B1(E[8]), .B2(n238), .ZN(n269) );
  NAND3_X1 U86 ( .A1(n271), .A2(n270), .A3(n269), .ZN(Y[8]) );
  AOI22_X1 U87 ( .A1(B[9]), .A2(n336), .B1(A[9]), .B2(n340), .ZN(n274) );
  NAND2_X1 U88 ( .A1(C[9]), .A2(n236), .ZN(n273) );
  AOI22_X1 U89 ( .A1(D[9]), .A2(n233), .B1(E[9]), .B2(n238), .ZN(n272) );
  NAND3_X1 U90 ( .A1(n274), .A2(n273), .A3(n272), .ZN(Y[9]) );
  AOI22_X1 U91 ( .A1(B[10]), .A2(n336), .B1(A[10]), .B2(n340), .ZN(n277) );
  NAND2_X1 U92 ( .A1(C[10]), .A2(n236), .ZN(n276) );
  AOI22_X1 U93 ( .A1(D[10]), .A2(n233), .B1(E[10]), .B2(n238), .ZN(n275) );
  NAND3_X1 U94 ( .A1(n277), .A2(n276), .A3(n275), .ZN(Y[10]) );
  AOI22_X1 U95 ( .A1(B[11]), .A2(n341), .B1(A[11]), .B2(n340), .ZN(n280) );
  NAND2_X1 U96 ( .A1(C[11]), .A2(n236), .ZN(n279) );
  AOI22_X1 U97 ( .A1(D[11]), .A2(n233), .B1(E[11]), .B2(n238), .ZN(n278) );
  NAND3_X1 U98 ( .A1(n280), .A2(n279), .A3(n278), .ZN(Y[11]) );
  AOI22_X1 U99 ( .A1(B[12]), .A2(n336), .B1(A[12]), .B2(n340), .ZN(n283) );
  NAND2_X1 U100 ( .A1(C[12]), .A2(n236), .ZN(n282) );
  AOI22_X1 U101 ( .A1(D[12]), .A2(n348), .B1(E[12]), .B2(n238), .ZN(n281) );
  AOI22_X1 U102 ( .A1(B[13]), .A2(n341), .B1(A[13]), .B2(n340), .ZN(n286) );
  NAND2_X1 U103 ( .A1(C[13]), .A2(n236), .ZN(n285) );
  AOI22_X1 U104 ( .A1(D[13]), .A2(n348), .B1(E[13]), .B2(n238), .ZN(n284) );
  NAND3_X1 U105 ( .A1(n286), .A2(n285), .A3(n284), .ZN(Y[13]) );
  AOI22_X1 U106 ( .A1(B[14]), .A2(n336), .B1(A[14]), .B2(n340), .ZN(n289) );
  NAND2_X1 U107 ( .A1(C[14]), .A2(n236), .ZN(n288) );
  AOI22_X1 U108 ( .A1(D[14]), .A2(n348), .B1(E[14]), .B2(n238), .ZN(n287) );
  NAND3_X1 U109 ( .A1(n289), .A2(n288), .A3(n287), .ZN(Y[14]) );
  AOI22_X1 U110 ( .A1(B[15]), .A2(n341), .B1(A[15]), .B2(n340), .ZN(n292) );
  AOI22_X1 U111 ( .A1(D[15]), .A2(n348), .B1(E[15]), .B2(n238), .ZN(n290) );
  NAND3_X1 U112 ( .A1(n292), .A2(n291), .A3(n290), .ZN(Y[15]) );
  NAND3_X1 U113 ( .A1(n295), .A2(n294), .A3(n293), .ZN(Y[16]) );
  AOI22_X1 U114 ( .A1(B[17]), .A2(n336), .B1(A[17]), .B2(n340), .ZN(n298) );
  NAND2_X1 U115 ( .A1(C[17]), .A2(n236), .ZN(n297) );
  AOI22_X1 U116 ( .A1(D[17]), .A2(n348), .B1(E[17]), .B2(n238), .ZN(n296) );
  NAND3_X1 U117 ( .A1(n298), .A2(n297), .A3(n296), .ZN(Y[17]) );
  AOI22_X1 U118 ( .A1(B[18]), .A2(n341), .B1(A[18]), .B2(n340), .ZN(n301) );
  NAND2_X1 U119 ( .A1(C[18]), .A2(n235), .ZN(n300) );
  AOI22_X1 U120 ( .A1(D[18]), .A2(n348), .B1(E[18]), .B2(n237), .ZN(n299) );
  NAND3_X1 U121 ( .A1(n301), .A2(n300), .A3(n299), .ZN(Y[18]) );
  AOI22_X1 U122 ( .A1(B[19]), .A2(n341), .B1(A[19]), .B2(n340), .ZN(n304) );
  NAND2_X1 U123 ( .A1(C[19]), .A2(n235), .ZN(n303) );
  AOI22_X1 U124 ( .A1(D[19]), .A2(n348), .B1(E[19]), .B2(n237), .ZN(n302) );
  NAND3_X1 U125 ( .A1(n304), .A2(n303), .A3(n302), .ZN(Y[19]) );
  AOI22_X1 U126 ( .A1(B[20]), .A2(n341), .B1(A[20]), .B2(n340), .ZN(n307) );
  NAND2_X1 U127 ( .A1(C[20]), .A2(n235), .ZN(n306) );
  AOI22_X1 U128 ( .A1(D[20]), .A2(n348), .B1(E[20]), .B2(n237), .ZN(n305) );
  NAND3_X1 U129 ( .A1(n307), .A2(n306), .A3(n305), .ZN(Y[20]) );
  AOI22_X1 U130 ( .A1(B[21]), .A2(n336), .B1(A[21]), .B2(n340), .ZN(n310) );
  NAND2_X1 U131 ( .A1(C[21]), .A2(n235), .ZN(n309) );
  AOI22_X1 U132 ( .A1(D[21]), .A2(n348), .B1(E[21]), .B2(n237), .ZN(n308) );
  NAND3_X1 U133 ( .A1(n310), .A2(n309), .A3(n308), .ZN(Y[21]) );
  AOI22_X1 U134 ( .A1(B[22]), .A2(n336), .B1(A[22]), .B2(n340), .ZN(n313) );
  NAND2_X1 U135 ( .A1(C[22]), .A2(n235), .ZN(n312) );
  AOI22_X1 U136 ( .A1(D[22]), .A2(n348), .B1(E[22]), .B2(n237), .ZN(n311) );
  NAND3_X1 U137 ( .A1(n313), .A2(n312), .A3(n311), .ZN(Y[22]) );
  AOI22_X1 U138 ( .A1(B[23]), .A2(n336), .B1(A[23]), .B2(n340), .ZN(n316) );
  NAND2_X1 U139 ( .A1(C[23]), .A2(n236), .ZN(n315) );
  AOI22_X1 U140 ( .A1(D[23]), .A2(n348), .B1(E[23]), .B2(n238), .ZN(n314) );
  NAND3_X1 U141 ( .A1(n316), .A2(n315), .A3(n314), .ZN(Y[23]) );
  AOI22_X1 U142 ( .A1(B[24]), .A2(n336), .B1(A[24]), .B2(n340), .ZN(n319) );
  AOI22_X1 U143 ( .A1(D[24]), .A2(n348), .B1(E[24]), .B2(n237), .ZN(n317) );
  NAND3_X1 U144 ( .A1(n319), .A2(n318), .A3(n317), .ZN(Y[24]) );
  NAND2_X1 U145 ( .A1(D[25]), .A2(n348), .ZN(n324) );
  INV_X1 U146 ( .A(A[25]), .ZN(n321) );
  OAI22_X1 U147 ( .A1(n346), .A2(n321), .B1(n345), .B2(n239), .ZN(n322) );
  AOI21_X1 U148 ( .B1(C[25]), .B2(n235), .A(n322), .ZN(n323) );
  NAND3_X1 U149 ( .A1(n325), .A2(n324), .A3(n323), .ZN(Y[25]) );
  NAND3_X1 U150 ( .A1(n328), .A2(n327), .A3(n326), .ZN(Y[26]) );
  NAND3_X1 U151 ( .A1(n332), .A2(n331), .A3(n330), .ZN(Y[27]) );
  NAND3_X1 U152 ( .A1(n339), .A2(n338), .A3(n337), .ZN(Y[29]) );
  NAND3_X1 U153 ( .A1(n344), .A2(n343), .A3(n342), .ZN(Y[30]) );
  NAND3_X1 U154 ( .A1(n351), .A2(n350), .A3(n349), .ZN(Y[31]) );
endmodule


module p4adder_N32_3 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  wire   [8:0] C;
  assign n1 = B[11];
  assign n2 = B[7];
  assign n3 = B[14];
  assign n4 = B[15];
  assign n5 = B[16];
  assign n6 = B[24];
  assign n7 = B[23];
  assign n8 = B[27];
  assign n9 = B[25];

  CarryGen_N32_3 Cgen ( .A(A), .B({B[31:29], n10, n8, B[26], n17, n18, n7, 
        B[22:17], n5, n4, n3, B[13:12], n1, B[10:8], n2, B[6:0]}), .Cin(Cin), 
        .C(C) );
  SumGen_N32_3 Sgen ( .A(A), .B({B[31:28], n20, B[26], n9, n6, n19, n13, 
        B[21:20], n15, B[18:17], n5, n16, n3, B[13:12], n14, B[10:8], n11, 
        B[6:4], n12, B[2:0]}), .C(C), .S(S), .Cout(Cout) );
  CLKBUF_X1 U1 ( .A(B[28]), .Z(n10) );
  CLKBUF_X1 U2 ( .A(n2), .Z(n11) );
  CLKBUF_X1 U3 ( .A(B[3]), .Z(n12) );
  BUF_X2 U4 ( .A(B[22]), .Z(n13) );
  CLKBUF_X1 U5 ( .A(n8), .Z(n20) );
  CLKBUF_X1 U6 ( .A(n1), .Z(n14) );
  BUF_X1 U7 ( .A(n9), .Z(n17) );
  CLKBUF_X1 U8 ( .A(B[19]), .Z(n15) );
  CLKBUF_X1 U9 ( .A(n4), .Z(n16) );
  CLKBUF_X1 U10 ( .A(n6), .Z(n18) );
  CLKBUF_X1 U11 ( .A(n7), .Z(n19) );
endmodule


module mux51_generic_N32_3 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351;

  INV_X2 U2 ( .A(n346), .ZN(n309) );
  NAND3_X2 U3 ( .A1(n324), .A2(n323), .A3(n322), .ZN(Y[25]) );
  BUF_X2 U4 ( .A(n222), .Z(n225) );
  BUF_X2 U5 ( .A(n348), .Z(n230) );
  BUF_X2 U6 ( .A(n344), .Z(n223) );
  BUF_X2 U7 ( .A(n348), .Z(n229) );
  BUF_X2 U8 ( .A(n222), .Z(n226) );
  NOR2_X1 U9 ( .A1(n346), .A2(n236), .ZN(n284) );
  BUF_X2 U10 ( .A(n344), .Z(n224) );
  NOR2_X1 U11 ( .A1(n346), .A2(n239), .ZN(n321) );
  NOR2_X1 U12 ( .A1(n346), .A2(n238), .ZN(n317) );
  NOR2_X1 U13 ( .A1(n346), .A2(n237), .ZN(n313) );
  NOR2_X1 U14 ( .A1(n346), .A2(n231), .ZN(n325) );
  NOR2_X1 U15 ( .A1(n346), .A2(n232), .ZN(n332) );
  NOR2_X1 U16 ( .A1(n346), .A2(n233), .ZN(n336) );
  NOR2_X1 U17 ( .A1(n346), .A2(n234), .ZN(n340) );
  NOR2_X1 U18 ( .A1(n346), .A2(n235), .ZN(n347) );
  NOR3_X1 U19 ( .A1(S[0]), .A2(n241), .A3(S[1]), .ZN(n348) );
  NOR3_X1 U20 ( .A1(S[0]), .A2(S[2]), .A3(S[1]), .ZN(n344) );
  NOR3_X1 U21 ( .A1(S[0]), .A2(S[2]), .A3(n240), .ZN(n345) );
  AND3_X1 U22 ( .A1(S[0]), .A2(n241), .A3(n240), .ZN(n222) );
  AOI21_X1 U23 ( .B1(E[29]), .B2(n229), .A(n336), .ZN(n337) );
  AOI21_X1 U24 ( .B1(E[31]), .B2(n229), .A(n347), .ZN(n349) );
  AOI21_X1 U25 ( .B1(E[30]), .B2(n229), .A(n340), .ZN(n341) );
  AOI21_X1 U26 ( .B1(E[14]), .B2(n229), .A(n284), .ZN(n285) );
  AOI21_X1 U27 ( .B1(E[28]), .B2(n229), .A(n332), .ZN(n333) );
  AOI22_X1 U28 ( .A1(A[27]), .A2(n223), .B1(B[27]), .B2(n225), .ZN(n329) );
  AOI22_X1 U29 ( .A1(D[27]), .A2(n309), .B1(E[27]), .B2(n229), .ZN(n331) );
  NAND2_X1 U30 ( .A1(C[27]), .A2(n227), .ZN(n330) );
  AOI21_X1 U31 ( .B1(E[23]), .B2(n229), .A(n313), .ZN(n314) );
  AOI21_X1 U32 ( .B1(E[26]), .B2(n229), .A(n325), .ZN(n326) );
  AOI21_X1 U33 ( .B1(E[25]), .B2(n229), .A(n321), .ZN(n322) );
  AOI21_X1 U34 ( .B1(E[24]), .B2(n229), .A(n317), .ZN(n318) );
  NAND3_X2 U35 ( .A1(S[0]), .A2(S[1]), .A3(n241), .ZN(n346) );
  CLKBUF_X3 U36 ( .A(n345), .Z(n227) );
  CLKBUF_X3 U37 ( .A(n345), .Z(n228) );
  INV_X1 U38 ( .A(D[26]), .ZN(n231) );
  INV_X1 U39 ( .A(D[28]), .ZN(n232) );
  INV_X1 U40 ( .A(D[29]), .ZN(n233) );
  INV_X1 U41 ( .A(D[30]), .ZN(n234) );
  INV_X1 U42 ( .A(D[31]), .ZN(n235) );
  INV_X1 U43 ( .A(D[14]), .ZN(n236) );
  INV_X1 U44 ( .A(D[23]), .ZN(n237) );
  INV_X1 U45 ( .A(D[24]), .ZN(n238) );
  INV_X1 U46 ( .A(D[25]), .ZN(n239) );
  INV_X1 U47 ( .A(S[2]), .ZN(n241) );
  INV_X1 U48 ( .A(S[1]), .ZN(n240) );
  AOI22_X1 U49 ( .A1(B[0]), .A2(n225), .B1(A[0]), .B2(n223), .ZN(n244) );
  NAND2_X1 U50 ( .A1(C[0]), .A2(n227), .ZN(n243) );
  AOI22_X1 U51 ( .A1(D[0]), .A2(n309), .B1(E[0]), .B2(n230), .ZN(n242) );
  NAND3_X1 U52 ( .A1(n244), .A2(n243), .A3(n242), .ZN(Y[0]) );
  AOI22_X1 U53 ( .A1(B[1]), .A2(n226), .B1(A[1]), .B2(n224), .ZN(n247) );
  NAND2_X1 U54 ( .A1(C[1]), .A2(n228), .ZN(n246) );
  AOI22_X1 U55 ( .A1(D[1]), .A2(n309), .B1(E[1]), .B2(n229), .ZN(n245) );
  NAND3_X1 U56 ( .A1(n247), .A2(n246), .A3(n245), .ZN(Y[1]) );
  AOI22_X1 U57 ( .A1(B[2]), .A2(n226), .B1(A[2]), .B2(n224), .ZN(n250) );
  NAND2_X1 U58 ( .A1(C[2]), .A2(n228), .ZN(n249) );
  AOI22_X1 U59 ( .A1(D[2]), .A2(n309), .B1(E[2]), .B2(n230), .ZN(n248) );
  NAND3_X1 U60 ( .A1(n250), .A2(n249), .A3(n248), .ZN(Y[2]) );
  AOI22_X1 U61 ( .A1(B[3]), .A2(n226), .B1(A[3]), .B2(n224), .ZN(n253) );
  NAND2_X1 U62 ( .A1(C[3]), .A2(n228), .ZN(n252) );
  AOI22_X1 U63 ( .A1(D[3]), .A2(n309), .B1(E[3]), .B2(n230), .ZN(n251) );
  NAND3_X1 U64 ( .A1(n253), .A2(n252), .A3(n251), .ZN(Y[3]) );
  AOI22_X1 U65 ( .A1(B[4]), .A2(n226), .B1(A[4]), .B2(n224), .ZN(n256) );
  NAND2_X1 U66 ( .A1(C[4]), .A2(n228), .ZN(n255) );
  AOI22_X1 U67 ( .A1(D[4]), .A2(n309), .B1(E[4]), .B2(n230), .ZN(n254) );
  NAND3_X1 U68 ( .A1(n256), .A2(n255), .A3(n254), .ZN(Y[4]) );
  AOI22_X1 U69 ( .A1(B[5]), .A2(n226), .B1(A[5]), .B2(n224), .ZN(n259) );
  NAND2_X1 U70 ( .A1(C[5]), .A2(n228), .ZN(n258) );
  AOI22_X1 U71 ( .A1(D[5]), .A2(n309), .B1(E[5]), .B2(n230), .ZN(n257) );
  NAND3_X1 U72 ( .A1(n259), .A2(n258), .A3(n257), .ZN(Y[5]) );
  AOI22_X1 U73 ( .A1(B[6]), .A2(n226), .B1(A[6]), .B2(n224), .ZN(n262) );
  NAND2_X1 U74 ( .A1(C[6]), .A2(n228), .ZN(n261) );
  AOI22_X1 U75 ( .A1(D[6]), .A2(n309), .B1(E[6]), .B2(n230), .ZN(n260) );
  NAND3_X1 U76 ( .A1(n262), .A2(n261), .A3(n260), .ZN(Y[6]) );
  AOI22_X1 U77 ( .A1(B[7]), .A2(n226), .B1(A[7]), .B2(n224), .ZN(n265) );
  NAND2_X1 U78 ( .A1(C[7]), .A2(n228), .ZN(n264) );
  AOI22_X1 U79 ( .A1(D[7]), .A2(n309), .B1(E[7]), .B2(n230), .ZN(n263) );
  NAND3_X1 U80 ( .A1(n265), .A2(n264), .A3(n263), .ZN(Y[7]) );
  AOI22_X1 U81 ( .A1(B[8]), .A2(n226), .B1(A[8]), .B2(n224), .ZN(n268) );
  NAND2_X1 U82 ( .A1(C[8]), .A2(n228), .ZN(n267) );
  AOI22_X1 U83 ( .A1(D[8]), .A2(n309), .B1(E[8]), .B2(n230), .ZN(n266) );
  NAND3_X1 U84 ( .A1(n268), .A2(n267), .A3(n266), .ZN(Y[8]) );
  AOI22_X1 U85 ( .A1(B[9]), .A2(n226), .B1(A[9]), .B2(n224), .ZN(n271) );
  NAND2_X1 U86 ( .A1(C[9]), .A2(n228), .ZN(n270) );
  AOI22_X1 U87 ( .A1(D[9]), .A2(n309), .B1(E[9]), .B2(n230), .ZN(n269) );
  NAND3_X1 U88 ( .A1(n271), .A2(n270), .A3(n269), .ZN(Y[9]) );
  AOI22_X1 U89 ( .A1(B[10]), .A2(n226), .B1(A[10]), .B2(n224), .ZN(n274) );
  NAND2_X1 U90 ( .A1(C[10]), .A2(n228), .ZN(n273) );
  AOI22_X1 U91 ( .A1(D[10]), .A2(n309), .B1(E[10]), .B2(n230), .ZN(n272) );
  NAND3_X1 U92 ( .A1(n274), .A2(n273), .A3(n272), .ZN(Y[10]) );
  AOI22_X1 U93 ( .A1(B[11]), .A2(n226), .B1(A[11]), .B2(n224), .ZN(n277) );
  NAND2_X1 U94 ( .A1(C[11]), .A2(n228), .ZN(n276) );
  AOI22_X1 U95 ( .A1(D[11]), .A2(n309), .B1(E[11]), .B2(n230), .ZN(n275) );
  NAND3_X1 U96 ( .A1(n277), .A2(n276), .A3(n275), .ZN(Y[11]) );
  AOI22_X1 U97 ( .A1(B[12]), .A2(n226), .B1(A[12]), .B2(n224), .ZN(n280) );
  NAND2_X1 U98 ( .A1(C[12]), .A2(n228), .ZN(n279) );
  AOI22_X1 U99 ( .A1(D[12]), .A2(n309), .B1(E[12]), .B2(n230), .ZN(n278) );
  NAND3_X1 U100 ( .A1(n280), .A2(n279), .A3(n278), .ZN(Y[12]) );
  AOI22_X1 U101 ( .A1(B[13]), .A2(n226), .B1(A[13]), .B2(n223), .ZN(n283) );
  NAND2_X1 U102 ( .A1(C[13]), .A2(n228), .ZN(n282) );
  AOI22_X1 U103 ( .A1(D[13]), .A2(n309), .B1(E[13]), .B2(n230), .ZN(n281) );
  NAND3_X1 U104 ( .A1(n283), .A2(n282), .A3(n281), .ZN(Y[13]) );
  AOI22_X1 U105 ( .A1(B[14]), .A2(n225), .B1(A[14]), .B2(n223), .ZN(n287) );
  NAND2_X1 U106 ( .A1(C[14]), .A2(n227), .ZN(n286) );
  NAND3_X1 U107 ( .A1(n287), .A2(n286), .A3(n285), .ZN(Y[14]) );
  AOI22_X1 U108 ( .A1(B[15]), .A2(n225), .B1(A[15]), .B2(n223), .ZN(n290) );
  NAND2_X1 U109 ( .A1(C[15]), .A2(n227), .ZN(n289) );
  AOI22_X1 U110 ( .A1(D[15]), .A2(n309), .B1(E[15]), .B2(n230), .ZN(n288) );
  NAND3_X1 U111 ( .A1(n290), .A2(n289), .A3(n288), .ZN(Y[15]) );
  AOI22_X1 U112 ( .A1(B[16]), .A2(n225), .B1(A[16]), .B2(n223), .ZN(n293) );
  NAND2_X1 U113 ( .A1(C[16]), .A2(n227), .ZN(n292) );
  AOI22_X1 U114 ( .A1(D[16]), .A2(n309), .B1(E[16]), .B2(n230), .ZN(n291) );
  NAND3_X1 U115 ( .A1(n293), .A2(n292), .A3(n291), .ZN(Y[16]) );
  AOI22_X1 U116 ( .A1(B[17]), .A2(n225), .B1(A[17]), .B2(n223), .ZN(n296) );
  NAND2_X1 U117 ( .A1(C[17]), .A2(n227), .ZN(n295) );
  AOI22_X1 U118 ( .A1(D[17]), .A2(n309), .B1(E[17]), .B2(n230), .ZN(n294) );
  NAND3_X1 U119 ( .A1(n296), .A2(n295), .A3(n294), .ZN(Y[17]) );
  AOI22_X1 U120 ( .A1(B[18]), .A2(n225), .B1(A[18]), .B2(n223), .ZN(n299) );
  NAND2_X1 U121 ( .A1(C[18]), .A2(n227), .ZN(n298) );
  AOI22_X1 U122 ( .A1(D[18]), .A2(n309), .B1(E[18]), .B2(n230), .ZN(n297) );
  NAND3_X1 U123 ( .A1(n299), .A2(n298), .A3(n297), .ZN(Y[18]) );
  AOI22_X1 U124 ( .A1(B[19]), .A2(n225), .B1(A[19]), .B2(n223), .ZN(n302) );
  NAND2_X1 U125 ( .A1(C[19]), .A2(n227), .ZN(n301) );
  AOI22_X1 U126 ( .A1(D[19]), .A2(n309), .B1(E[19]), .B2(n230), .ZN(n300) );
  NAND3_X1 U127 ( .A1(n302), .A2(n301), .A3(n300), .ZN(Y[19]) );
  AOI22_X1 U128 ( .A1(B[20]), .A2(n225), .B1(A[20]), .B2(n223), .ZN(n305) );
  NAND2_X1 U129 ( .A1(C[20]), .A2(n227), .ZN(n304) );
  AOI22_X1 U130 ( .A1(D[20]), .A2(n309), .B1(E[20]), .B2(n230), .ZN(n303) );
  NAND3_X1 U131 ( .A1(n305), .A2(n304), .A3(n303), .ZN(Y[20]) );
  AOI22_X1 U132 ( .A1(B[21]), .A2(n225), .B1(A[21]), .B2(n223), .ZN(n308) );
  NAND2_X1 U133 ( .A1(C[21]), .A2(n227), .ZN(n307) );
  AOI22_X1 U134 ( .A1(D[21]), .A2(n309), .B1(E[21]), .B2(n229), .ZN(n306) );
  NAND3_X1 U135 ( .A1(n308), .A2(n307), .A3(n306), .ZN(Y[21]) );
  AOI22_X1 U136 ( .A1(B[22]), .A2(n225), .B1(A[22]), .B2(n223), .ZN(n312) );
  NAND2_X1 U137 ( .A1(C[22]), .A2(n227), .ZN(n311) );
  AOI22_X1 U138 ( .A1(D[22]), .A2(n309), .B1(E[22]), .B2(n229), .ZN(n310) );
  NAND3_X1 U139 ( .A1(n312), .A2(n311), .A3(n310), .ZN(Y[22]) );
  AOI22_X1 U140 ( .A1(B[23]), .A2(n225), .B1(A[23]), .B2(n223), .ZN(n316) );
  NAND2_X1 U141 ( .A1(C[23]), .A2(n227), .ZN(n315) );
  NAND3_X1 U142 ( .A1(n316), .A2(n315), .A3(n314), .ZN(Y[23]) );
  AOI22_X1 U143 ( .A1(B[24]), .A2(n225), .B1(A[24]), .B2(n223), .ZN(n320) );
  NAND2_X1 U144 ( .A1(C[24]), .A2(n227), .ZN(n319) );
  NAND3_X1 U145 ( .A1(n320), .A2(n319), .A3(n318), .ZN(Y[24]) );
  AOI22_X1 U146 ( .A1(B[25]), .A2(n225), .B1(A[25]), .B2(n223), .ZN(n324) );
  NAND2_X1 U147 ( .A1(C[25]), .A2(n227), .ZN(n323) );
  AOI22_X1 U148 ( .A1(B[26]), .A2(n225), .B1(A[26]), .B2(n223), .ZN(n328) );
  NAND2_X1 U149 ( .A1(C[26]), .A2(n227), .ZN(n327) );
  NAND3_X1 U150 ( .A1(n328), .A2(n327), .A3(n326), .ZN(Y[26]) );
  NAND3_X1 U151 ( .A1(n331), .A2(n330), .A3(n329), .ZN(Y[27]) );
  AOI22_X1 U152 ( .A1(B[28]), .A2(n225), .B1(A[28]), .B2(n223), .ZN(n335) );
  NAND2_X1 U153 ( .A1(C[28]), .A2(n227), .ZN(n334) );
  NAND3_X1 U154 ( .A1(n335), .A2(n334), .A3(n333), .ZN(Y[28]) );
  AOI22_X1 U155 ( .A1(B[29]), .A2(n225), .B1(A[29]), .B2(n223), .ZN(n339) );
  NAND2_X1 U156 ( .A1(C[29]), .A2(n227), .ZN(n338) );
  NAND3_X1 U157 ( .A1(n339), .A2(n338), .A3(n337), .ZN(Y[29]) );
  AOI22_X1 U158 ( .A1(B[30]), .A2(n225), .B1(A[30]), .B2(n223), .ZN(n343) );
  NAND2_X1 U159 ( .A1(C[30]), .A2(n227), .ZN(n342) );
  NAND3_X1 U160 ( .A1(n343), .A2(n342), .A3(n341), .ZN(Y[30]) );
  AOI22_X1 U161 ( .A1(B[31]), .A2(n225), .B1(A[31]), .B2(n223), .ZN(n351) );
  NAND2_X1 U162 ( .A1(C[31]), .A2(n227), .ZN(n350) );
  NAND3_X1 U163 ( .A1(n351), .A2(n350), .A3(n349), .ZN(Y[31]) );
endmodule


module p4adder_N32_4 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  wire   [8:0] C;
  assign n1 = B[27];
  assign n2 = B[12];
  assign n3 = B[15];
  assign n5 = B[7];
  assign n6 = B[20];
  assign n7 = B[16];
  assign n8 = B[11];
  assign n9 = B[24];
  assign n10 = B[23];
  assign n11 = B[19];

  CarryGen_N32_4 Cgen ( .A(A), .B({B[31:28], n1, B[26:25], n17, n10, B[22:21], 
        n6, n11, B[18:17], n7, n3, B[14:13], n2, n8, B[10:8], n5, B[6:0]}), 
        .Cin(Cin), .C(C) );
  SumGen_N32_4 Sgen ( .A(A), .B({B[31:28], n13, B[26:25], n9, n15, B[22:21], 
        n6, n20, B[18:17], n7, n19, n14, B[13], n2, n18, B[10:8], n16, B[6:4], 
        n12, B[2:0]}), .C(C), .S(S), .Cout(Cout) );
  CLKBUF_X1 U1 ( .A(n1), .Z(n13) );
  CLKBUF_X1 U2 ( .A(B[3]), .Z(n12) );
  BUF_X1 U3 ( .A(n9), .Z(n17) );
  BUF_X1 U4 ( .A(B[14]), .Z(n14) );
  CLKBUF_X1 U5 ( .A(n10), .Z(n15) );
  CLKBUF_X1 U6 ( .A(n5), .Z(n16) );
  CLKBUF_X1 U7 ( .A(n8), .Z(n18) );
  CLKBUF_X1 U8 ( .A(n3), .Z(n19) );
  CLKBUF_X1 U9 ( .A(n11), .Z(n20) );
endmodule


module mux51_generic_N32_4 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419;

  INV_X2 U2 ( .A(n349), .ZN(n416) );
  BUF_X2 U3 ( .A(n225), .Z(n232) );
  NAND3_X2 U4 ( .A1(n365), .A2(n364), .A3(n363), .ZN(Y[21]) );
  NAND3_X2 U5 ( .A1(n286), .A2(n285), .A3(n284), .ZN(Y[8]) );
  CLKBUF_X1 U6 ( .A(n225), .Z(n233) );
  BUF_X2 U7 ( .A(n416), .Z(n235) );
  NAND2_X1 U8 ( .A1(C[11]), .A2(n235), .ZN(n297) );
  BUF_X2 U9 ( .A(n411), .Z(n231) );
  NOR2_X1 U10 ( .A1(n349), .A2(n327), .ZN(n330) );
  NAND2_X1 U11 ( .A1(n258), .A2(n257), .ZN(n414) );
  CLKBUF_X1 U12 ( .A(n411), .Z(n229) );
  BUF_X1 U13 ( .A(n411), .Z(n230) );
  NOR2_X1 U14 ( .A1(n349), .A2(n299), .ZN(n302) );
  NOR2_X1 U15 ( .A1(n349), .A2(n306), .ZN(n309) );
  NOR2_X1 U16 ( .A1(n349), .A2(n313), .ZN(n316) );
  CLKBUF_X1 U17 ( .A(n225), .Z(n234) );
  NOR3_X1 U18 ( .A1(S[0]), .A2(n259), .A3(S[1]), .ZN(n411) );
  AND3_X1 U19 ( .A1(S[0]), .A2(S[1]), .A3(n259), .ZN(n225) );
  AOI21_X1 U20 ( .B1(C[29]), .B2(n416), .A(n402), .ZN(n403) );
  AOI21_X1 U21 ( .B1(C[25]), .B2(n416), .A(n382), .ZN(n383) );
  AOI21_X1 U22 ( .B1(C[26]), .B2(n416), .A(n387), .ZN(n388) );
  AOI21_X1 U23 ( .B1(C[27]), .B2(n416), .A(n392), .ZN(n393) );
  AOI21_X1 U24 ( .B1(C[28]), .B2(n416), .A(n397), .ZN(n398) );
  AOI21_X1 U25 ( .B1(C[30]), .B2(n416), .A(n407), .ZN(n408) );
  AOI21_X1 U26 ( .B1(C[31]), .B2(n416), .A(n415), .ZN(n417) );
  AOI21_X1 U27 ( .B1(C[24]), .B2(n416), .A(n377), .ZN(n378) );
  AOI21_X1 U28 ( .B1(C[20]), .B2(n235), .A(n357), .ZN(n358) );
  AOI21_X1 U29 ( .B1(C[23]), .B2(n416), .A(n372), .ZN(n373) );
  AOI21_X1 U30 ( .B1(C[22]), .B2(n416), .A(n367), .ZN(n368) );
  NAND3_X1 U31 ( .A1(S[0]), .A2(n259), .A3(n256), .ZN(n226) );
  NAND3_X1 U32 ( .A1(S[0]), .A2(n259), .A3(n256), .ZN(n227) );
  NAND2_X2 U33 ( .A1(n258), .A2(n257), .ZN(n228) );
  NAND3_X2 U34 ( .A1(S[1]), .A2(n259), .A3(n258), .ZN(n349) );
  INV_X1 U35 ( .A(B[15]), .ZN(n236) );
  INV_X1 U36 ( .A(B[14]), .ZN(n237) );
  INV_X1 U37 ( .A(B[23]), .ZN(n238) );
  INV_X1 U38 ( .A(B[24]), .ZN(n239) );
  INV_X1 U39 ( .A(B[25]), .ZN(n240) );
  INV_X1 U40 ( .A(B[26]), .ZN(n241) );
  INV_X1 U41 ( .A(B[27]), .ZN(n242) );
  INV_X1 U42 ( .A(B[28]), .ZN(n243) );
  INV_X1 U43 ( .A(B[29]), .ZN(n244) );
  INV_X1 U44 ( .A(B[30]), .ZN(n245) );
  INV_X1 U45 ( .A(B[31]), .ZN(n246) );
  INV_X1 U46 ( .A(B[12]), .ZN(n247) );
  INV_X1 U47 ( .A(B[13]), .ZN(n248) );
  INV_X1 U48 ( .A(B[16]), .ZN(n249) );
  INV_X1 U49 ( .A(B[17]), .ZN(n250) );
  INV_X1 U50 ( .A(B[18]), .ZN(n251) );
  INV_X1 U51 ( .A(B[19]), .ZN(n252) );
  INV_X1 U52 ( .A(B[20]), .ZN(n253) );
  INV_X1 U53 ( .A(B[21]), .ZN(n254) );
  INV_X1 U54 ( .A(B[22]), .ZN(n255) );
  INV_X1 U55 ( .A(S[2]), .ZN(n259) );
  INV_X1 U56 ( .A(S[1]), .ZN(n256) );
  NAND3_X1 U57 ( .A1(S[0]), .A2(n259), .A3(n256), .ZN(n412) );
  INV_X1 U58 ( .A(n412), .ZN(n294) );
  INV_X1 U59 ( .A(S[0]), .ZN(n258) );
  NOR2_X1 U60 ( .A1(S[2]), .A2(S[1]), .ZN(n257) );
  INV_X1 U61 ( .A(n228), .ZN(n293) );
  AOI22_X1 U62 ( .A1(B[0]), .A2(n294), .B1(A[0]), .B2(n293), .ZN(n262) );
  NAND2_X1 U63 ( .A1(C[0]), .A2(n235), .ZN(n261) );
  AOI22_X1 U64 ( .A1(D[0]), .A2(n232), .B1(E[0]), .B2(n231), .ZN(n260) );
  NAND3_X1 U65 ( .A1(n262), .A2(n261), .A3(n260), .ZN(Y[0]) );
  AOI22_X1 U66 ( .A1(B[1]), .A2(n294), .B1(A[1]), .B2(n293), .ZN(n265) );
  NAND2_X1 U67 ( .A1(C[1]), .A2(n235), .ZN(n264) );
  AOI22_X1 U68 ( .A1(D[1]), .A2(n232), .B1(E[1]), .B2(n231), .ZN(n263) );
  NAND3_X1 U69 ( .A1(n265), .A2(n264), .A3(n263), .ZN(Y[1]) );
  AOI22_X1 U70 ( .A1(B[2]), .A2(n294), .B1(A[2]), .B2(n293), .ZN(n268) );
  NAND2_X1 U71 ( .A1(C[2]), .A2(n235), .ZN(n267) );
  AOI22_X1 U72 ( .A1(D[2]), .A2(n232), .B1(E[2]), .B2(n231), .ZN(n266) );
  NAND3_X1 U73 ( .A1(n268), .A2(n267), .A3(n266), .ZN(Y[2]) );
  AOI22_X1 U74 ( .A1(B[3]), .A2(n294), .B1(A[3]), .B2(n293), .ZN(n271) );
  NAND2_X1 U75 ( .A1(C[3]), .A2(n235), .ZN(n270) );
  AOI22_X1 U76 ( .A1(D[3]), .A2(n232), .B1(E[3]), .B2(n231), .ZN(n269) );
  NAND3_X1 U77 ( .A1(n271), .A2(n270), .A3(n269), .ZN(Y[3]) );
  AOI22_X1 U78 ( .A1(B[4]), .A2(n294), .B1(A[4]), .B2(n293), .ZN(n274) );
  NAND2_X1 U79 ( .A1(C[4]), .A2(n235), .ZN(n273) );
  AOI22_X1 U80 ( .A1(D[4]), .A2(n232), .B1(E[4]), .B2(n231), .ZN(n272) );
  NAND3_X1 U81 ( .A1(n274), .A2(n273), .A3(n272), .ZN(Y[4]) );
  AOI22_X1 U82 ( .A1(B[5]), .A2(n294), .B1(A[5]), .B2(n293), .ZN(n277) );
  NAND2_X1 U83 ( .A1(C[5]), .A2(n235), .ZN(n276) );
  AOI22_X1 U84 ( .A1(D[5]), .A2(n232), .B1(E[5]), .B2(n231), .ZN(n275) );
  NAND3_X1 U85 ( .A1(n277), .A2(n276), .A3(n275), .ZN(Y[5]) );
  AOI22_X1 U86 ( .A1(B[6]), .A2(n294), .B1(A[6]), .B2(n293), .ZN(n280) );
  NAND2_X1 U87 ( .A1(C[6]), .A2(n235), .ZN(n279) );
  AOI22_X1 U88 ( .A1(D[6]), .A2(n232), .B1(E[6]), .B2(n231), .ZN(n278) );
  NAND3_X1 U89 ( .A1(n280), .A2(n279), .A3(n278), .ZN(Y[6]) );
  AOI22_X1 U90 ( .A1(B[7]), .A2(n294), .B1(A[7]), .B2(n293), .ZN(n283) );
  NAND2_X1 U91 ( .A1(C[7]), .A2(n235), .ZN(n282) );
  AOI22_X1 U92 ( .A1(D[7]), .A2(n232), .B1(E[7]), .B2(n231), .ZN(n281) );
  NAND3_X1 U93 ( .A1(n283), .A2(n282), .A3(n281), .ZN(Y[7]) );
  AOI22_X1 U94 ( .A1(B[8]), .A2(n294), .B1(A[8]), .B2(n293), .ZN(n286) );
  NAND2_X1 U95 ( .A1(C[8]), .A2(n235), .ZN(n285) );
  AOI22_X1 U96 ( .A1(D[8]), .A2(n232), .B1(E[8]), .B2(n230), .ZN(n284) );
  AOI22_X1 U97 ( .A1(B[9]), .A2(n294), .B1(A[9]), .B2(n293), .ZN(n289) );
  NAND2_X1 U98 ( .A1(C[9]), .A2(n235), .ZN(n288) );
  AOI22_X1 U99 ( .A1(D[9]), .A2(n232), .B1(E[9]), .B2(n230), .ZN(n287) );
  NAND3_X1 U100 ( .A1(n289), .A2(n288), .A3(n287), .ZN(Y[9]) );
  AOI22_X1 U101 ( .A1(B[10]), .A2(n294), .B1(A[10]), .B2(n293), .ZN(n292) );
  NAND2_X1 U102 ( .A1(C[10]), .A2(n235), .ZN(n291) );
  AOI22_X1 U103 ( .A1(D[10]), .A2(n232), .B1(E[10]), .B2(n230), .ZN(n290) );
  NAND3_X1 U104 ( .A1(n292), .A2(n291), .A3(n290), .ZN(Y[10]) );
  AOI22_X1 U105 ( .A1(B[11]), .A2(n294), .B1(A[11]), .B2(n293), .ZN(n298) );
  NAND2_X1 U106 ( .A1(E[11]), .A2(n230), .ZN(n296) );
  NAND2_X1 U107 ( .A1(D[11]), .A2(n232), .ZN(n295) );
  NAND4_X1 U108 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[11]) );
  NAND2_X1 U109 ( .A1(E[12]), .A2(n230), .ZN(n305) );
  NAND2_X1 U110 ( .A1(D[12]), .A2(n233), .ZN(n304) );
  INV_X1 U111 ( .A(C[12]), .ZN(n299) );
  INV_X1 U112 ( .A(A[12]), .ZN(n300) );
  OAI22_X1 U113 ( .A1(n228), .A2(n300), .B1(n226), .B2(n247), .ZN(n301) );
  NOR2_X1 U114 ( .A1(n302), .A2(n301), .ZN(n303) );
  NAND3_X1 U115 ( .A1(n305), .A2(n304), .A3(n303), .ZN(Y[12]) );
  NAND2_X1 U116 ( .A1(E[13]), .A2(n230), .ZN(n312) );
  NAND2_X1 U117 ( .A1(D[13]), .A2(n233), .ZN(n311) );
  INV_X1 U118 ( .A(C[13]), .ZN(n306) );
  INV_X1 U119 ( .A(A[13]), .ZN(n307) );
  OAI22_X1 U120 ( .A1(n414), .A2(n307), .B1(n227), .B2(n248), .ZN(n308) );
  NOR2_X1 U121 ( .A1(n309), .A2(n308), .ZN(n310) );
  NAND3_X1 U122 ( .A1(n312), .A2(n311), .A3(n310), .ZN(Y[13]) );
  NAND2_X1 U123 ( .A1(E[14]), .A2(n230), .ZN(n319) );
  NAND2_X1 U124 ( .A1(D[14]), .A2(n233), .ZN(n318) );
  INV_X1 U125 ( .A(C[14]), .ZN(n313) );
  INV_X1 U126 ( .A(A[14]), .ZN(n314) );
  OAI22_X1 U127 ( .A1(n228), .A2(n314), .B1(n412), .B2(n237), .ZN(n315) );
  NOR2_X1 U128 ( .A1(n316), .A2(n315), .ZN(n317) );
  NAND3_X1 U129 ( .A1(n319), .A2(n318), .A3(n317), .ZN(Y[14]) );
  NAND2_X1 U130 ( .A1(E[15]), .A2(n230), .ZN(n326) );
  NAND2_X1 U131 ( .A1(D[15]), .A2(n233), .ZN(n325) );
  INV_X1 U132 ( .A(C[15]), .ZN(n320) );
  NOR2_X1 U133 ( .A1(n349), .A2(n320), .ZN(n323) );
  INV_X1 U134 ( .A(A[15]), .ZN(n321) );
  OAI22_X1 U135 ( .A1(n414), .A2(n321), .B1(n226), .B2(n236), .ZN(n322) );
  NOR2_X1 U136 ( .A1(n323), .A2(n322), .ZN(n324) );
  NAND3_X1 U137 ( .A1(n326), .A2(n325), .A3(n324), .ZN(Y[15]) );
  NAND2_X1 U138 ( .A1(E[16]), .A2(n230), .ZN(n333) );
  NAND2_X1 U139 ( .A1(D[16]), .A2(n233), .ZN(n332) );
  INV_X1 U140 ( .A(C[16]), .ZN(n327) );
  INV_X1 U141 ( .A(A[16]), .ZN(n328) );
  OAI22_X1 U142 ( .A1(n228), .A2(n328), .B1(n227), .B2(n249), .ZN(n329) );
  NOR2_X1 U143 ( .A1(n330), .A2(n329), .ZN(n331) );
  NAND3_X1 U144 ( .A1(n333), .A2(n332), .A3(n331), .ZN(Y[16]) );
  NAND2_X1 U145 ( .A1(E[17]), .A2(n230), .ZN(n340) );
  NAND2_X1 U146 ( .A1(D[17]), .A2(n233), .ZN(n339) );
  INV_X1 U147 ( .A(C[17]), .ZN(n334) );
  NOR2_X1 U148 ( .A1(n349), .A2(n334), .ZN(n337) );
  INV_X1 U149 ( .A(A[17]), .ZN(n335) );
  OAI22_X1 U150 ( .A1(n414), .A2(n335), .B1(n412), .B2(n250), .ZN(n336) );
  NOR2_X1 U151 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND3_X1 U152 ( .A1(n340), .A2(n339), .A3(n338), .ZN(Y[17]) );
  NAND2_X1 U153 ( .A1(E[18]), .A2(n230), .ZN(n347) );
  NAND2_X1 U154 ( .A1(D[18]), .A2(n233), .ZN(n346) );
  INV_X1 U155 ( .A(C[18]), .ZN(n341) );
  NOR2_X1 U156 ( .A1(n349), .A2(n341), .ZN(n344) );
  INV_X1 U157 ( .A(A[18]), .ZN(n342) );
  OAI22_X1 U158 ( .A1(n228), .A2(n342), .B1(n226), .B2(n251), .ZN(n343) );
  NOR2_X1 U159 ( .A1(n344), .A2(n343), .ZN(n345) );
  NAND3_X1 U160 ( .A1(n347), .A2(n346), .A3(n345), .ZN(Y[18]) );
  NAND2_X1 U161 ( .A1(E[19]), .A2(n230), .ZN(n355) );
  NAND2_X1 U162 ( .A1(D[19]), .A2(n233), .ZN(n354) );
  INV_X1 U163 ( .A(C[19]), .ZN(n348) );
  NOR2_X1 U164 ( .A1(n349), .A2(n348), .ZN(n352) );
  INV_X1 U165 ( .A(A[19]), .ZN(n350) );
  OAI22_X1 U166 ( .A1(n414), .A2(n350), .B1(n227), .B2(n252), .ZN(n351) );
  NOR2_X1 U167 ( .A1(n352), .A2(n351), .ZN(n353) );
  NAND3_X1 U168 ( .A1(n355), .A2(n354), .A3(n353), .ZN(Y[19]) );
  NAND2_X1 U169 ( .A1(E[20]), .A2(n229), .ZN(n360) );
  NAND2_X1 U170 ( .A1(D[20]), .A2(n233), .ZN(n359) );
  INV_X1 U171 ( .A(A[20]), .ZN(n356) );
  OAI22_X1 U172 ( .A1(n228), .A2(n356), .B1(n412), .B2(n253), .ZN(n357) );
  NAND3_X1 U173 ( .A1(n360), .A2(n359), .A3(n358), .ZN(Y[20]) );
  NAND2_X1 U174 ( .A1(E[21]), .A2(n229), .ZN(n365) );
  NAND2_X1 U175 ( .A1(D[21]), .A2(n233), .ZN(n364) );
  INV_X1 U176 ( .A(A[21]), .ZN(n361) );
  OAI22_X1 U177 ( .A1(n414), .A2(n361), .B1(n226), .B2(n254), .ZN(n362) );
  AOI21_X1 U178 ( .B1(C[21]), .B2(n235), .A(n362), .ZN(n363) );
  NAND2_X1 U179 ( .A1(E[22]), .A2(n229), .ZN(n370) );
  NAND2_X1 U180 ( .A1(D[22]), .A2(n233), .ZN(n369) );
  INV_X1 U181 ( .A(A[22]), .ZN(n366) );
  OAI22_X1 U182 ( .A1(n228), .A2(n366), .B1(n227), .B2(n255), .ZN(n367) );
  NAND3_X1 U183 ( .A1(n370), .A2(n369), .A3(n368), .ZN(Y[22]) );
  NAND2_X1 U184 ( .A1(E[23]), .A2(n229), .ZN(n375) );
  NAND2_X1 U185 ( .A1(D[23]), .A2(n233), .ZN(n374) );
  INV_X1 U186 ( .A(A[23]), .ZN(n371) );
  OAI22_X1 U187 ( .A1(n414), .A2(n371), .B1(n412), .B2(n238), .ZN(n372) );
  NAND3_X1 U188 ( .A1(n375), .A2(n374), .A3(n373), .ZN(Y[23]) );
  NAND2_X1 U189 ( .A1(E[24]), .A2(n229), .ZN(n380) );
  NAND2_X1 U190 ( .A1(D[24]), .A2(n234), .ZN(n379) );
  INV_X1 U191 ( .A(A[24]), .ZN(n376) );
  OAI22_X1 U192 ( .A1(n228), .A2(n376), .B1(n226), .B2(n239), .ZN(n377) );
  NAND3_X1 U193 ( .A1(n380), .A2(n379), .A3(n378), .ZN(Y[24]) );
  NAND2_X1 U194 ( .A1(E[25]), .A2(n229), .ZN(n385) );
  NAND2_X1 U195 ( .A1(D[25]), .A2(n234), .ZN(n384) );
  INV_X1 U196 ( .A(A[25]), .ZN(n381) );
  OAI22_X1 U197 ( .A1(n414), .A2(n381), .B1(n227), .B2(n240), .ZN(n382) );
  NAND3_X1 U198 ( .A1(n385), .A2(n384), .A3(n383), .ZN(Y[25]) );
  NAND2_X1 U199 ( .A1(E[26]), .A2(n229), .ZN(n390) );
  NAND2_X1 U200 ( .A1(D[26]), .A2(n234), .ZN(n389) );
  INV_X1 U201 ( .A(A[26]), .ZN(n386) );
  OAI22_X1 U202 ( .A1(n228), .A2(n386), .B1(n412), .B2(n241), .ZN(n387) );
  NAND3_X1 U203 ( .A1(n390), .A2(n389), .A3(n388), .ZN(Y[26]) );
  NAND2_X1 U204 ( .A1(E[27]), .A2(n229), .ZN(n395) );
  NAND2_X1 U205 ( .A1(D[27]), .A2(n234), .ZN(n394) );
  INV_X1 U206 ( .A(A[27]), .ZN(n391) );
  OAI22_X1 U207 ( .A1(n414), .A2(n391), .B1(n226), .B2(n242), .ZN(n392) );
  NAND3_X1 U208 ( .A1(n395), .A2(n394), .A3(n393), .ZN(Y[27]) );
  NAND2_X1 U209 ( .A1(E[28]), .A2(n229), .ZN(n400) );
  NAND2_X1 U210 ( .A1(D[28]), .A2(n234), .ZN(n399) );
  INV_X1 U211 ( .A(A[28]), .ZN(n396) );
  OAI22_X1 U212 ( .A1(n228), .A2(n396), .B1(n227), .B2(n243), .ZN(n397) );
  NAND3_X1 U213 ( .A1(n400), .A2(n399), .A3(n398), .ZN(Y[28]) );
  NAND2_X1 U214 ( .A1(E[29]), .A2(n229), .ZN(n405) );
  NAND2_X1 U215 ( .A1(D[29]), .A2(n234), .ZN(n404) );
  INV_X1 U216 ( .A(A[29]), .ZN(n401) );
  OAI22_X1 U217 ( .A1(n414), .A2(n401), .B1(n412), .B2(n244), .ZN(n402) );
  NAND3_X1 U218 ( .A1(n405), .A2(n404), .A3(n403), .ZN(Y[29]) );
  NAND2_X1 U219 ( .A1(E[30]), .A2(n229), .ZN(n410) );
  NAND2_X1 U220 ( .A1(D[30]), .A2(n234), .ZN(n409) );
  INV_X1 U221 ( .A(A[30]), .ZN(n406) );
  OAI22_X1 U222 ( .A1(n228), .A2(n406), .B1(n226), .B2(n245), .ZN(n407) );
  NAND3_X1 U223 ( .A1(n410), .A2(n409), .A3(n408), .ZN(Y[30]) );
  NAND2_X1 U224 ( .A1(E[31]), .A2(n229), .ZN(n419) );
  NAND2_X1 U225 ( .A1(D[31]), .A2(n234), .ZN(n418) );
  INV_X1 U226 ( .A(A[31]), .ZN(n413) );
  OAI22_X1 U227 ( .A1(n414), .A2(n413), .B1(n227), .B2(n246), .ZN(n415) );
  NAND3_X1 U228 ( .A1(n419), .A2(n418), .A3(n417), .ZN(Y[31]) );
endmodule


module p4adder_N32_5 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [8:0] C;
  assign n1 = B[4];
  assign n2 = B[16];
  assign n3 = B[3];
  assign n4 = B[23];
  assign n5 = B[7];
  assign n6 = B[11];
  assign n7 = B[19];
  assign n8 = B[15];

  CarryGen_N32_5 Cgen ( .A(A), .B({B[31:24], n4, B[22:20], n7, B[18:17], n17, 
        n8, B[14:12], n6, B[10:8], n5, B[6:5], n11, n3, B[2], n9, B[0]}), 
        .Cin(Cin), .C(C) );
  SumGen_N32_5 Sgen ( .A(A), .B({B[31:24], n16, B[22:20], n13, B[18:17], n2, 
        n18, n14, B[13:12], n19, B[10:8], n12, n15, B[5], n1, n10, B[2:0]}), 
        .C(C), .S(S), .Cout(Cout) );
  CLKBUF_X1 U1 ( .A(B[1]), .Z(n9) );
  BUF_X2 U2 ( .A(B[6]), .Z(n15) );
  BUF_X1 U3 ( .A(n3), .Z(n10) );
  CLKBUF_X1 U4 ( .A(n1), .Z(n11) );
  CLKBUF_X1 U5 ( .A(n5), .Z(n12) );
  CLKBUF_X1 U6 ( .A(n4), .Z(n16) );
  CLKBUF_X1 U7 ( .A(n7), .Z(n13) );
  CLKBUF_X1 U8 ( .A(n2), .Z(n17) );
  BUF_X2 U9 ( .A(B[14]), .Z(n14) );
  CLKBUF_X1 U10 ( .A(n8), .Z(n18) );
  CLKBUF_X1 U11 ( .A(n6), .Z(n19) );
endmodule


module mux51_generic_N32_5 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418;

  BUF_X1 U2 ( .A(n233), .Z(n236) );
  NAND4_X2 U3 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .ZN(Y[4]) );
  NAND4_X2 U4 ( .A1(n304), .A2(n303), .A3(n302), .A4(n301), .ZN(Y[8]) );
  BUF_X1 U5 ( .A(n414), .Z(n234) );
  BUF_X2 U6 ( .A(n414), .Z(n235) );
  AND2_X1 U7 ( .A1(E[18]), .A2(n237), .ZN(n232) );
  BUF_X2 U8 ( .A(n233), .Z(n237) );
  NOR2_X1 U9 ( .A1(n415), .A2(n258), .ZN(n314) );
  NOR2_X1 U10 ( .A1(n415), .A2(n240), .ZN(n377) );
  NOR2_X1 U11 ( .A1(n415), .A2(n241), .ZN(n382) );
  NOR2_X1 U12 ( .A1(n415), .A2(n239), .ZN(n372) );
  NOR2_X1 U13 ( .A1(n415), .A2(n244), .ZN(n397) );
  NOR2_X1 U14 ( .A1(n415), .A2(n243), .ZN(n392) );
  NOR2_X1 U15 ( .A1(n415), .A2(n242), .ZN(n387) );
  NOR2_X1 U16 ( .A1(n415), .A2(n245), .ZN(n402) );
  NOR2_X1 U17 ( .A1(n415), .A2(n246), .ZN(n407) );
  NOR2_X1 U18 ( .A1(n415), .A2(n247), .ZN(n416) );
  NOR2_X1 U19 ( .A1(n415), .A2(n260), .ZN(n345) );
  NOR2_X1 U20 ( .A1(n415), .A2(n263), .ZN(n361) );
  NOR2_X1 U21 ( .A1(n415), .A2(n238), .ZN(n367) );
  NOR2_X1 U22 ( .A1(n415), .A2(n261), .ZN(n355) );
  AND2_X1 U23 ( .A1(n268), .A2(n267), .ZN(n233) );
  AOI21_X1 U24 ( .B1(E[10]), .B2(n236), .A(n314), .ZN(n315) );
  NOR2_X1 U25 ( .A1(n310), .A2(n309), .ZN(n313) );
  AOI21_X1 U26 ( .B1(C[22]), .B2(n234), .A(n366), .ZN(n369) );
  AOI21_X1 U27 ( .B1(C[28]), .B2(n234), .A(n396), .ZN(n399) );
  AOI21_X1 U28 ( .B1(E[28]), .B2(n236), .A(n397), .ZN(n398) );
  AOI21_X1 U29 ( .B1(C[29]), .B2(n234), .A(n401), .ZN(n404) );
  AOI21_X1 U30 ( .B1(E[29]), .B2(n236), .A(n402), .ZN(n403) );
  AOI21_X1 U31 ( .B1(C[30]), .B2(n234), .A(n406), .ZN(n409) );
  AOI21_X1 U32 ( .B1(E[30]), .B2(n236), .A(n407), .ZN(n408) );
  AOI21_X1 U33 ( .B1(C[31]), .B2(n234), .A(n413), .ZN(n418) );
  AOI21_X1 U34 ( .B1(E[31]), .B2(n236), .A(n416), .ZN(n417) );
  AOI21_X1 U35 ( .B1(C[24]), .B2(n234), .A(n376), .ZN(n379) );
  AOI21_X1 U36 ( .B1(E[24]), .B2(n236), .A(n377), .ZN(n378) );
  AOI21_X1 U37 ( .B1(C[27]), .B2(n234), .A(n391), .ZN(n394) );
  AOI21_X1 U38 ( .B1(E[27]), .B2(n236), .A(n392), .ZN(n393) );
  AOI21_X1 U39 ( .B1(C[23]), .B2(n234), .A(n371), .ZN(n374) );
  AOI21_X1 U40 ( .B1(E[23]), .B2(n236), .A(n372), .ZN(n373) );
  AOI21_X1 U41 ( .B1(C[25]), .B2(n234), .A(n381), .ZN(n384) );
  AOI21_X1 U42 ( .B1(E[25]), .B2(n236), .A(n382), .ZN(n383) );
  AOI21_X1 U43 ( .B1(C[26]), .B2(n234), .A(n386), .ZN(n389) );
  AOI21_X1 U44 ( .B1(E[26]), .B2(n236), .A(n387), .ZN(n388) );
  NAND2_X1 U45 ( .A1(C[9]), .A2(n234), .ZN(n307) );
  NAND4_X1 U46 ( .A1(n340), .A2(n339), .A3(n338), .A4(n337), .ZN(Y[16]) );
  NAND2_X1 U47 ( .A1(E[19]), .A2(n237), .ZN(n353) );
  NAND2_X1 U48 ( .A1(C[18]), .A2(n235), .ZN(n347) );
  AOI21_X1 U49 ( .B1(E[22]), .B2(n236), .A(n367), .ZN(n368) );
  NAND2_X1 U50 ( .A1(C[21]), .A2(n235), .ZN(n363) );
  NAND2_X1 U51 ( .A1(C[20]), .A2(n234), .ZN(n357) );
  AOI21_X1 U52 ( .B1(E[21]), .B2(n237), .A(n361), .ZN(n362) );
  AOI21_X1 U53 ( .B1(E[20]), .B2(n236), .A(n355), .ZN(n356) );
  NAND3_X2 U54 ( .A1(S[0]), .A2(n266), .A3(n264), .ZN(n410) );
  NAND3_X2 U55 ( .A1(S[0]), .A2(S[1]), .A3(n266), .ZN(n415) );
  INV_X1 U56 ( .A(D[22]), .ZN(n238) );
  INV_X1 U57 ( .A(D[23]), .ZN(n239) );
  INV_X1 U58 ( .A(D[24]), .ZN(n240) );
  INV_X1 U59 ( .A(D[25]), .ZN(n241) );
  INV_X1 U60 ( .A(D[26]), .ZN(n242) );
  INV_X1 U61 ( .A(D[27]), .ZN(n243) );
  INV_X1 U62 ( .A(D[28]), .ZN(n244) );
  INV_X1 U63 ( .A(D[29]), .ZN(n245) );
  INV_X1 U64 ( .A(D[30]), .ZN(n246) );
  INV_X1 U65 ( .A(D[31]), .ZN(n247) );
  INV_X1 U66 ( .A(B[22]), .ZN(n248) );
  INV_X1 U67 ( .A(B[23]), .ZN(n249) );
  INV_X1 U68 ( .A(B[24]), .ZN(n250) );
  INV_X1 U69 ( .A(B[25]), .ZN(n251) );
  INV_X1 U70 ( .A(B[26]), .ZN(n252) );
  INV_X1 U71 ( .A(B[27]), .ZN(n253) );
  INV_X1 U72 ( .A(B[28]), .ZN(n254) );
  INV_X1 U73 ( .A(B[29]), .ZN(n255) );
  INV_X1 U74 ( .A(B[30]), .ZN(n256) );
  INV_X1 U75 ( .A(B[31]), .ZN(n257) );
  INV_X1 U76 ( .A(D[10]), .ZN(n258) );
  INV_X1 U77 ( .A(B[10]), .ZN(n259) );
  INV_X1 U78 ( .A(D[18]), .ZN(n260) );
  INV_X1 U79 ( .A(D[20]), .ZN(n261) );
  INV_X1 U80 ( .A(B[19]), .ZN(n262) );
  INV_X1 U81 ( .A(D[21]), .ZN(n263) );
  INV_X1 U82 ( .A(S[2]), .ZN(n266) );
  INV_X1 U83 ( .A(S[1]), .ZN(n264) );
  INV_X1 U84 ( .A(n410), .ZN(n360) );
  INV_X1 U85 ( .A(S[0]), .ZN(n268) );
  NOR2_X1 U86 ( .A1(S[2]), .A2(S[1]), .ZN(n265) );
  NAND2_X2 U87 ( .A1(n268), .A2(n265), .ZN(n412) );
  INV_X1 U88 ( .A(n412), .ZN(n359) );
  AOI22_X1 U89 ( .A1(B[0]), .A2(n360), .B1(A[0]), .B2(n359), .ZN(n272) );
  NAND3_X1 U90 ( .A1(S[1]), .A2(n266), .A3(n268), .ZN(n310) );
  INV_X1 U91 ( .A(n310), .ZN(n414) );
  NAND2_X1 U92 ( .A1(C[0]), .A2(n235), .ZN(n271) );
  INV_X1 U93 ( .A(n415), .ZN(n349) );
  NAND2_X1 U94 ( .A1(D[0]), .A2(n349), .ZN(n270) );
  NOR2_X1 U95 ( .A1(n266), .A2(S[1]), .ZN(n267) );
  NAND2_X1 U96 ( .A1(E[0]), .A2(n237), .ZN(n269) );
  NAND4_X1 U97 ( .A1(n272), .A2(n271), .A3(n270), .A4(n269), .ZN(Y[0]) );
  AOI22_X1 U98 ( .A1(B[1]), .A2(n360), .B1(A[1]), .B2(n359), .ZN(n276) );
  NAND2_X1 U99 ( .A1(C[1]), .A2(n235), .ZN(n275) );
  NAND2_X1 U100 ( .A1(D[1]), .A2(n349), .ZN(n274) );
  NAND2_X1 U101 ( .A1(E[1]), .A2(n237), .ZN(n273) );
  NAND4_X1 U102 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .ZN(Y[1]) );
  AOI22_X1 U103 ( .A1(B[2]), .A2(n360), .B1(A[2]), .B2(n359), .ZN(n280) );
  NAND2_X1 U104 ( .A1(C[2]), .A2(n235), .ZN(n279) );
  NAND2_X1 U105 ( .A1(D[2]), .A2(n349), .ZN(n278) );
  NAND2_X1 U106 ( .A1(E[2]), .A2(n236), .ZN(n277) );
  NAND4_X1 U107 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .ZN(Y[2]) );
  AOI22_X1 U108 ( .A1(B[3]), .A2(n360), .B1(A[3]), .B2(n359), .ZN(n284) );
  NAND2_X1 U109 ( .A1(C[3]), .A2(n235), .ZN(n283) );
  NAND2_X1 U110 ( .A1(D[3]), .A2(n349), .ZN(n282) );
  NAND2_X1 U111 ( .A1(E[3]), .A2(n237), .ZN(n281) );
  NAND4_X1 U112 ( .A1(n284), .A2(n283), .A3(n282), .A4(n281), .ZN(Y[3]) );
  AOI22_X1 U113 ( .A1(B[4]), .A2(n360), .B1(A[4]), .B2(n359), .ZN(n288) );
  NAND2_X1 U114 ( .A1(C[4]), .A2(n235), .ZN(n287) );
  NAND2_X1 U115 ( .A1(D[4]), .A2(n349), .ZN(n286) );
  NAND2_X1 U116 ( .A1(E[4]), .A2(n237), .ZN(n285) );
  AOI22_X1 U117 ( .A1(B[5]), .A2(n360), .B1(A[5]), .B2(n359), .ZN(n292) );
  NAND2_X1 U118 ( .A1(C[5]), .A2(n235), .ZN(n291) );
  NAND2_X1 U119 ( .A1(D[5]), .A2(n349), .ZN(n290) );
  NAND2_X1 U120 ( .A1(E[5]), .A2(n237), .ZN(n289) );
  NAND4_X1 U121 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(Y[5]) );
  AOI22_X1 U122 ( .A1(B[6]), .A2(n360), .B1(A[6]), .B2(n359), .ZN(n296) );
  NAND2_X1 U123 ( .A1(C[6]), .A2(n235), .ZN(n295) );
  NAND2_X1 U124 ( .A1(D[6]), .A2(n349), .ZN(n294) );
  NAND2_X1 U125 ( .A1(E[6]), .A2(n237), .ZN(n293) );
  NAND4_X1 U126 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(Y[6]) );
  AOI22_X1 U127 ( .A1(B[7]), .A2(n360), .B1(A[7]), .B2(n359), .ZN(n300) );
  NAND2_X1 U128 ( .A1(C[7]), .A2(n235), .ZN(n299) );
  NAND2_X1 U129 ( .A1(D[7]), .A2(n349), .ZN(n298) );
  NAND2_X1 U130 ( .A1(E[7]), .A2(n237), .ZN(n297) );
  NAND4_X1 U131 ( .A1(n300), .A2(n299), .A3(n298), .A4(n297), .ZN(Y[7]) );
  AOI22_X1 U132 ( .A1(B[8]), .A2(n360), .B1(A[8]), .B2(n359), .ZN(n304) );
  NAND2_X1 U133 ( .A1(C[8]), .A2(n235), .ZN(n303) );
  NAND2_X1 U134 ( .A1(D[8]), .A2(n349), .ZN(n302) );
  NAND2_X1 U135 ( .A1(E[8]), .A2(n237), .ZN(n301) );
  AOI22_X1 U136 ( .A1(B[9]), .A2(n360), .B1(A[9]), .B2(n359), .ZN(n308) );
  NAND2_X1 U137 ( .A1(D[9]), .A2(n349), .ZN(n306) );
  NAND2_X1 U138 ( .A1(E[9]), .A2(n237), .ZN(n305) );
  NAND4_X1 U139 ( .A1(n308), .A2(n307), .A3(n306), .A4(n305), .ZN(Y[9]) );
  INV_X1 U140 ( .A(C[10]), .ZN(n309) );
  INV_X1 U141 ( .A(A[10]), .ZN(n311) );
  OAI22_X1 U142 ( .A1(n412), .A2(n311), .B1(n410), .B2(n259), .ZN(n312) );
  NOR2_X1 U143 ( .A1(n313), .A2(n312), .ZN(n316) );
  NAND2_X1 U144 ( .A1(n316), .A2(n315), .ZN(Y[10]) );
  AOI22_X1 U145 ( .A1(B[11]), .A2(n360), .B1(A[11]), .B2(n359), .ZN(n320) );
  NAND2_X1 U146 ( .A1(C[11]), .A2(n235), .ZN(n319) );
  NAND2_X1 U147 ( .A1(D[11]), .A2(n349), .ZN(n318) );
  NAND2_X1 U148 ( .A1(E[11]), .A2(n237), .ZN(n317) );
  NAND4_X1 U149 ( .A1(n320), .A2(n319), .A3(n318), .A4(n317), .ZN(Y[11]) );
  AOI22_X1 U150 ( .A1(B[12]), .A2(n360), .B1(A[12]), .B2(n359), .ZN(n324) );
  NAND2_X1 U151 ( .A1(C[12]), .A2(n235), .ZN(n323) );
  NAND2_X1 U152 ( .A1(D[12]), .A2(n349), .ZN(n322) );
  NAND2_X1 U153 ( .A1(E[12]), .A2(n237), .ZN(n321) );
  NAND4_X1 U154 ( .A1(n324), .A2(n323), .A3(n322), .A4(n321), .ZN(Y[12]) );
  AOI22_X1 U155 ( .A1(B[13]), .A2(n360), .B1(A[13]), .B2(n359), .ZN(n328) );
  NAND2_X1 U156 ( .A1(C[13]), .A2(n235), .ZN(n327) );
  NAND2_X1 U157 ( .A1(D[13]), .A2(n349), .ZN(n326) );
  NAND2_X1 U158 ( .A1(E[13]), .A2(n237), .ZN(n325) );
  NAND4_X1 U159 ( .A1(n328), .A2(n327), .A3(n326), .A4(n325), .ZN(Y[13]) );
  AOI22_X1 U160 ( .A1(B[14]), .A2(n360), .B1(A[14]), .B2(n359), .ZN(n332) );
  NAND2_X1 U161 ( .A1(C[14]), .A2(n235), .ZN(n331) );
  NAND2_X1 U162 ( .A1(D[14]), .A2(n349), .ZN(n330) );
  NAND2_X1 U163 ( .A1(E[14]), .A2(n237), .ZN(n329) );
  NAND4_X1 U164 ( .A1(n332), .A2(n331), .A3(n330), .A4(n329), .ZN(Y[14]) );
  AOI22_X1 U165 ( .A1(B[15]), .A2(n360), .B1(A[15]), .B2(n359), .ZN(n336) );
  NAND2_X1 U166 ( .A1(C[15]), .A2(n235), .ZN(n335) );
  NAND2_X1 U167 ( .A1(D[15]), .A2(n349), .ZN(n334) );
  NAND2_X1 U168 ( .A1(E[15]), .A2(n237), .ZN(n333) );
  NAND4_X1 U169 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .ZN(Y[15]) );
  AOI22_X1 U170 ( .A1(B[16]), .A2(n360), .B1(A[16]), .B2(n359), .ZN(n340) );
  NAND2_X1 U171 ( .A1(C[16]), .A2(n235), .ZN(n339) );
  NAND2_X1 U172 ( .A1(D[16]), .A2(n349), .ZN(n338) );
  NAND2_X1 U173 ( .A1(E[16]), .A2(n237), .ZN(n337) );
  AOI22_X1 U174 ( .A1(B[17]), .A2(n360), .B1(A[17]), .B2(n359), .ZN(n344) );
  NAND2_X1 U175 ( .A1(C[17]), .A2(n235), .ZN(n343) );
  NAND2_X1 U176 ( .A1(D[17]), .A2(n349), .ZN(n342) );
  NAND2_X1 U177 ( .A1(E[17]), .A2(n237), .ZN(n341) );
  NAND4_X1 U178 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .ZN(Y[17]) );
  AOI22_X1 U179 ( .A1(B[18]), .A2(n360), .B1(A[18]), .B2(n359), .ZN(n348) );
  NOR2_X1 U180 ( .A1(n232), .A2(n345), .ZN(n346) );
  NAND3_X1 U181 ( .A1(n348), .A2(n347), .A3(n346), .ZN(Y[18]) );
  NAND2_X1 U182 ( .A1(D[19]), .A2(n349), .ZN(n354) );
  INV_X1 U183 ( .A(A[19]), .ZN(n350) );
  OAI22_X1 U184 ( .A1(n412), .A2(n350), .B1(n410), .B2(n262), .ZN(n351) );
  AOI21_X1 U185 ( .B1(C[19]), .B2(n235), .A(n351), .ZN(n352) );
  NAND3_X1 U186 ( .A1(n354), .A2(n353), .A3(n352), .ZN(Y[19]) );
  AOI22_X1 U187 ( .A1(B[20]), .A2(n360), .B1(A[20]), .B2(n359), .ZN(n358) );
  NAND3_X1 U188 ( .A1(n358), .A2(n357), .A3(n356), .ZN(Y[20]) );
  AOI22_X1 U189 ( .A1(B[21]), .A2(n360), .B1(A[21]), .B2(n359), .ZN(n364) );
  NAND3_X1 U190 ( .A1(n364), .A2(n363), .A3(n362), .ZN(Y[21]) );
  INV_X1 U191 ( .A(A[22]), .ZN(n365) );
  OAI22_X1 U192 ( .A1(n412), .A2(n365), .B1(n410), .B2(n248), .ZN(n366) );
  NAND2_X1 U193 ( .A1(n369), .A2(n368), .ZN(Y[22]) );
  INV_X1 U194 ( .A(A[23]), .ZN(n370) );
  OAI22_X1 U195 ( .A1(n412), .A2(n370), .B1(n410), .B2(n249), .ZN(n371) );
  NAND2_X1 U196 ( .A1(n374), .A2(n373), .ZN(Y[23]) );
  INV_X1 U197 ( .A(A[24]), .ZN(n375) );
  OAI22_X1 U198 ( .A1(n412), .A2(n375), .B1(n410), .B2(n250), .ZN(n376) );
  NAND2_X1 U199 ( .A1(n379), .A2(n378), .ZN(Y[24]) );
  INV_X1 U200 ( .A(A[25]), .ZN(n380) );
  OAI22_X1 U201 ( .A1(n412), .A2(n380), .B1(n410), .B2(n251), .ZN(n381) );
  NAND2_X1 U202 ( .A1(n384), .A2(n383), .ZN(Y[25]) );
  INV_X1 U203 ( .A(A[26]), .ZN(n385) );
  OAI22_X1 U204 ( .A1(n412), .A2(n385), .B1(n410), .B2(n252), .ZN(n386) );
  NAND2_X1 U205 ( .A1(n389), .A2(n388), .ZN(Y[26]) );
  INV_X1 U206 ( .A(A[27]), .ZN(n390) );
  OAI22_X1 U207 ( .A1(n412), .A2(n390), .B1(n410), .B2(n253), .ZN(n391) );
  NAND2_X1 U208 ( .A1(n394), .A2(n393), .ZN(Y[27]) );
  INV_X1 U209 ( .A(A[28]), .ZN(n395) );
  OAI22_X1 U210 ( .A1(n412), .A2(n395), .B1(n410), .B2(n254), .ZN(n396) );
  NAND2_X1 U211 ( .A1(n399), .A2(n398), .ZN(Y[28]) );
  INV_X1 U212 ( .A(A[29]), .ZN(n400) );
  OAI22_X1 U213 ( .A1(n412), .A2(n400), .B1(n410), .B2(n255), .ZN(n401) );
  NAND2_X1 U214 ( .A1(n404), .A2(n403), .ZN(Y[29]) );
  INV_X1 U215 ( .A(A[30]), .ZN(n405) );
  OAI22_X1 U216 ( .A1(n412), .A2(n405), .B1(n410), .B2(n256), .ZN(n406) );
  NAND2_X1 U217 ( .A1(n409), .A2(n408), .ZN(Y[30]) );
  INV_X1 U218 ( .A(A[31]), .ZN(n411) );
  OAI22_X1 U219 ( .A1(n412), .A2(n411), .B1(n410), .B2(n257), .ZN(n413) );
  NAND2_X1 U220 ( .A1(n418), .A2(n417), .ZN(Y[31]) );
endmodule


module Boothencoder_5 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   n9, n10, n11;

  OAI21_X1 U1 ( .B1(B[0]), .B2(B[1]), .A(n11), .ZN(n10) );
  NAND2_X1 U2 ( .A1(B[1]), .A2(B[0]), .ZN(n11) );
  AND3_X1 U3 ( .A1(n11), .A2(B[2]), .A3(n10), .ZN(S[2]) );
  AOI21_X1 U4 ( .B1(n11), .B2(n10), .A(B[2]), .ZN(S[0]) );
  MUX2_X1 U5 ( .A(n11), .B(n10), .S(B[2]), .Z(n9) );
  INV_X1 U6 ( .A(n9), .ZN(S[1]) );
endmodule


module p4adder_N32_6 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;
  wire   [8:0] C;
  assign n1 = B[8];
  assign n2 = A[0];
  assign n3 = B[11];
  assign n4 = B[0];
  assign n5 = B[7];
  assign n6 = B[15];
  assign n7 = B[3];

  CarryGen_N32_6 Cgen ( .A({A[31:1], n9}), .B({B[31:16], n6, B[14:12], n3, 
        B[10:9], n10, n5, B[6:4], n7, B[2:1], n8}), .Cin(Cin), .C(C) );
  SumGen_N32_6 Sgen ( .A({A[31:1], n2}), .B({B[31:16], n13, n11, B[13:12], n3, 
        B[10:9], n1, n14, B[6:4], n12, B[2:1], n4}), .C(C), .S(S), .Cout(Cout)
         );
  CLKBUF_X1 U1 ( .A(n4), .Z(n8) );
  CLKBUF_X1 U2 ( .A(n2), .Z(n9) );
  CLKBUF_X1 U3 ( .A(n7), .Z(n12) );
  CLKBUF_X1 U4 ( .A(n1), .Z(n10) );
  BUF_X1 U5 ( .A(B[14]), .Z(n11) );
  CLKBUF_X1 U6 ( .A(n6), .Z(n13) );
  CLKBUF_X1 U7 ( .A(n5), .Z(n14) );
endmodule


module mux51_generic_N32_6 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496;

  AND3_X2 U2 ( .A1(S[0]), .A2(n311), .A3(n312), .ZN(n241) );
  INV_X2 U3 ( .A(n241), .ZN(n252) );
  INV_X2 U4 ( .A(n491), .ZN(n239) );
  AND3_X2 U5 ( .A1(S[2]), .A2(n311), .A3(n310), .ZN(n243) );
  BUF_X4 U6 ( .A(n243), .Z(n245) );
  AND2_X1 U7 ( .A1(n310), .A2(n308), .ZN(n242) );
  NAND3_X2 U8 ( .A1(n343), .A2(n342), .A3(n341), .ZN(Y[4]) );
  NAND3_X2 U9 ( .A1(n429), .A2(n428), .A3(n427), .ZN(Y[20]) );
  BUF_X4 U10 ( .A(n242), .Z(n247) );
  INV_X1 U11 ( .A(n491), .ZN(n396) );
  NAND2_X4 U12 ( .A1(n309), .A2(n310), .ZN(n491) );
  NOR2_X1 U13 ( .A1(n249), .A2(n282), .ZN(n345) );
  NOR2_X1 U14 ( .A1(n249), .A2(n288), .ZN(n360) );
  NOR2_X1 U15 ( .A1(n251), .A2(n283), .ZN(n339) );
  NOR2_X1 U16 ( .A1(n251), .A2(n289), .ZN(n354) );
  NOR2_X1 U17 ( .A1(n251), .A2(n295), .ZN(n379) );
  NOR2_X1 U18 ( .A1(n250), .A2(n294), .ZN(n385) );
  CLKBUF_X1 U19 ( .A(n242), .Z(n246) );
  BUF_X2 U20 ( .A(n243), .Z(n244) );
  NOR2_X1 U21 ( .A1(n249), .A2(n286), .ZN(n355) );
  NOR2_X1 U22 ( .A1(n249), .A2(n290), .ZN(n365) );
  NOR2_X1 U23 ( .A1(n249), .A2(n292), .ZN(n370) );
  NOR2_X1 U24 ( .A1(n249), .A2(n255), .ZN(n375) );
  NOR2_X1 U25 ( .A1(n249), .A2(n253), .ZN(n380) );
  NOR2_X1 U26 ( .A1(n251), .A2(n287), .ZN(n349) );
  NOR2_X1 U27 ( .A1(n251), .A2(n293), .ZN(n364) );
  NOR2_X1 U28 ( .A1(n251), .A2(n256), .ZN(n369) );
  NOR2_X1 U29 ( .A1(n251), .A2(n291), .ZN(n359) );
  NOR2_X1 U30 ( .A1(n251), .A2(n254), .ZN(n374) );
  NOR2_X1 U31 ( .A1(n250), .A2(n298), .ZN(n395) );
  NOR2_X1 U32 ( .A1(n250), .A2(n296), .ZN(n390) );
  NOR2_X1 U33 ( .A1(n252), .A2(n297), .ZN(n384) );
  NOR2_X1 U34 ( .A1(n252), .A2(n301), .ZN(n394) );
  NOR2_X1 U35 ( .A1(n252), .A2(n299), .ZN(n389) );
  CLKBUF_X1 U36 ( .A(n242), .Z(n248) );
  AND3_X1 U37 ( .A1(S[0]), .A2(S[1]), .A3(n312), .ZN(n240) );
  NOR2_X1 U38 ( .A1(n249), .A2(n284), .ZN(n350) );
  NOR2_X1 U39 ( .A1(n251), .A2(n285), .ZN(n344) );
  NAND2_X1 U40 ( .A1(E[24]), .A2(n244), .ZN(n453) );
  NAND2_X1 U41 ( .A1(C[24]), .A2(n246), .ZN(n452) );
  NAND2_X1 U42 ( .A1(E[25]), .A2(n244), .ZN(n459) );
  NAND2_X1 U43 ( .A1(C[25]), .A2(n246), .ZN(n458) );
  NAND2_X1 U44 ( .A1(E[21]), .A2(n244), .ZN(n435) );
  NAND2_X1 U45 ( .A1(C[21]), .A2(n246), .ZN(n434) );
  NAND2_X1 U46 ( .A1(E[23]), .A2(n244), .ZN(n447) );
  NAND2_X1 U47 ( .A1(C[23]), .A2(n246), .ZN(n446) );
  NAND2_X1 U48 ( .A1(E[22]), .A2(n245), .ZN(n441) );
  NAND2_X1 U49 ( .A1(C[22]), .A2(n246), .ZN(n440) );
  NAND2_X1 U50 ( .A1(E[27]), .A2(n244), .ZN(n471) );
  NAND2_X1 U51 ( .A1(C[27]), .A2(n246), .ZN(n470) );
  NAND2_X1 U52 ( .A1(E[26]), .A2(n244), .ZN(n465) );
  NAND2_X1 U53 ( .A1(C[26]), .A2(n246), .ZN(n464) );
  NAND2_X1 U54 ( .A1(C[20]), .A2(n246), .ZN(n428) );
  NAND2_X1 U55 ( .A1(E[28]), .A2(n244), .ZN(n477) );
  NAND2_X1 U56 ( .A1(C[28]), .A2(n246), .ZN(n476) );
  NAND2_X1 U57 ( .A1(E[29]), .A2(n244), .ZN(n483) );
  NAND2_X1 U58 ( .A1(C[29]), .A2(n246), .ZN(n482) );
  NAND2_X1 U59 ( .A1(E[30]), .A2(n244), .ZN(n489) );
  NAND2_X1 U60 ( .A1(C[30]), .A2(n246), .ZN(n488) );
  NAND2_X1 U61 ( .A1(E[31]), .A2(n244), .ZN(n496) );
  NAND2_X1 U62 ( .A1(C[31]), .A2(n246), .ZN(n495) );
  NAND2_X1 U63 ( .A1(D[0]), .A2(n240), .ZN(n313) );
  NAND2_X1 U64 ( .A1(B[0]), .A2(n241), .ZN(n314) );
  AOI22_X1 U65 ( .A1(E[0]), .A2(n244), .B1(C[0]), .B2(n247), .ZN(n316) );
  NOR2_X1 U66 ( .A1(n491), .A2(n412), .ZN(n414) );
  NOR2_X1 U67 ( .A1(n491), .A2(n418), .ZN(n420) );
  NOR2_X1 U68 ( .A1(n491), .A2(n406), .ZN(n408) );
  NOR2_X1 U69 ( .A1(n491), .A2(n400), .ZN(n402) );
  NOR2_X1 U70 ( .A1(n491), .A2(n448), .ZN(n450) );
  NOR2_X1 U71 ( .A1(n491), .A2(n454), .ZN(n456) );
  NOR2_X1 U72 ( .A1(n491), .A2(n442), .ZN(n444) );
  NOR2_X1 U73 ( .A1(n491), .A2(n436), .ZN(n438) );
  NOR2_X1 U74 ( .A1(n491), .A2(n430), .ZN(n432) );
  NOR2_X1 U75 ( .A1(n491), .A2(n424), .ZN(n426) );
  NAND2_X1 U76 ( .A1(A[0]), .A2(n396), .ZN(n315) );
  NOR2_X1 U77 ( .A1(n249), .A2(n338), .ZN(n340) );
  NOR2_X1 U78 ( .A1(n249), .A2(n317), .ZN(n320) );
  NOR2_X1 U79 ( .A1(n249), .A2(n324), .ZN(n327) );
  NOR2_X1 U80 ( .A1(n249), .A2(n331), .ZN(n334) );
  NOR2_X1 U81 ( .A1(n251), .A2(n318), .ZN(n319) );
  NOR2_X1 U82 ( .A1(n251), .A2(n325), .ZN(n326) );
  NOR2_X1 U83 ( .A1(n251), .A2(n332), .ZN(n333) );
  NOR2_X1 U84 ( .A1(n491), .A2(n472), .ZN(n474) );
  NOR2_X1 U85 ( .A1(n491), .A2(n460), .ZN(n462) );
  NOR2_X1 U86 ( .A1(n491), .A2(n466), .ZN(n468) );
  NOR2_X1 U87 ( .A1(n491), .A2(n478), .ZN(n480) );
  NOR2_X1 U88 ( .A1(n491), .A2(n484), .ZN(n486) );
  NOR2_X1 U89 ( .A1(n491), .A2(n490), .ZN(n493) );
  NAND2_X1 U90 ( .A1(C[16]), .A2(n247), .ZN(n404) );
  NAND2_X1 U91 ( .A1(E[17]), .A2(n245), .ZN(n411) );
  NAND2_X1 U92 ( .A1(E[20]), .A2(n244), .ZN(n429) );
  NAND2_X1 U93 ( .A1(C[19]), .A2(n247), .ZN(n422) );
  NAND2_X1 U94 ( .A1(E[19]), .A2(n245), .ZN(n423) );
  NAND2_X1 U95 ( .A1(C[18]), .A2(n247), .ZN(n416) );
  INV_X2 U96 ( .A(n240), .ZN(n249) );
  INV_X2 U97 ( .A(n240), .ZN(n250) );
  INV_X2 U98 ( .A(n241), .ZN(n251) );
  INV_X1 U99 ( .A(D[12]), .ZN(n253) );
  INV_X1 U100 ( .A(B[11]), .ZN(n254) );
  INV_X1 U101 ( .A(D[11]), .ZN(n255) );
  INV_X1 U102 ( .A(B[10]), .ZN(n256) );
  INV_X1 U103 ( .A(D[20]), .ZN(n257) );
  INV_X1 U104 ( .A(D[21]), .ZN(n258) );
  INV_X1 U105 ( .A(D[22]), .ZN(n259) );
  INV_X1 U106 ( .A(D[23]), .ZN(n260) );
  INV_X1 U107 ( .A(D[24]), .ZN(n261) );
  INV_X1 U108 ( .A(D[25]), .ZN(n262) );
  INV_X1 U109 ( .A(D[26]), .ZN(n263) );
  INV_X1 U110 ( .A(D[27]), .ZN(n264) );
  INV_X1 U111 ( .A(D[28]), .ZN(n265) );
  INV_X1 U112 ( .A(D[29]), .ZN(n266) );
  INV_X1 U113 ( .A(D[30]), .ZN(n267) );
  INV_X1 U114 ( .A(D[31]), .ZN(n268) );
  INV_X1 U115 ( .A(B[19]), .ZN(n269) );
  INV_X1 U116 ( .A(B[20]), .ZN(n270) );
  INV_X1 U117 ( .A(B[21]), .ZN(n271) );
  INV_X1 U118 ( .A(B[22]), .ZN(n272) );
  INV_X1 U119 ( .A(B[23]), .ZN(n273) );
  INV_X1 U120 ( .A(B[24]), .ZN(n274) );
  INV_X1 U121 ( .A(B[25]), .ZN(n275) );
  INV_X1 U122 ( .A(B[26]), .ZN(n276) );
  INV_X1 U123 ( .A(B[27]), .ZN(n277) );
  INV_X1 U124 ( .A(B[28]), .ZN(n278) );
  INV_X1 U125 ( .A(B[29]), .ZN(n279) );
  INV_X1 U126 ( .A(B[30]), .ZN(n280) );
  INV_X1 U127 ( .A(B[31]), .ZN(n281) );
  INV_X1 U128 ( .A(D[5]), .ZN(n282) );
  INV_X1 U129 ( .A(B[4]), .ZN(n283) );
  INV_X1 U130 ( .A(D[6]), .ZN(n284) );
  INV_X1 U131 ( .A(B[5]), .ZN(n285) );
  INV_X1 U132 ( .A(D[7]), .ZN(n286) );
  INV_X1 U133 ( .A(B[6]), .ZN(n287) );
  INV_X1 U134 ( .A(D[8]), .ZN(n288) );
  INV_X1 U135 ( .A(B[7]), .ZN(n289) );
  INV_X1 U136 ( .A(D[9]), .ZN(n290) );
  INV_X1 U137 ( .A(B[8]), .ZN(n291) );
  INV_X1 U138 ( .A(D[10]), .ZN(n292) );
  INV_X1 U139 ( .A(B[9]), .ZN(n293) );
  INV_X1 U140 ( .A(D[13]), .ZN(n294) );
  INV_X1 U141 ( .A(B[12]), .ZN(n295) );
  INV_X1 U142 ( .A(D[14]), .ZN(n296) );
  INV_X1 U143 ( .A(B[13]), .ZN(n297) );
  INV_X1 U144 ( .A(D[15]), .ZN(n298) );
  INV_X1 U145 ( .A(B[14]), .ZN(n299) );
  INV_X1 U146 ( .A(D[16]), .ZN(n300) );
  INV_X1 U147 ( .A(B[15]), .ZN(n301) );
  INV_X1 U148 ( .A(D[17]), .ZN(n302) );
  INV_X1 U149 ( .A(B[16]), .ZN(n303) );
  INV_X1 U150 ( .A(D[18]), .ZN(n304) );
  INV_X1 U151 ( .A(B[17]), .ZN(n305) );
  INV_X1 U152 ( .A(D[19]), .ZN(n306) );
  INV_X1 U153 ( .A(B[18]), .ZN(n307) );
  INV_X1 U154 ( .A(S[1]), .ZN(n311) );
  INV_X1 U155 ( .A(S[0]), .ZN(n310) );
  NOR2_X1 U156 ( .A1(n311), .A2(S[2]), .ZN(n308) );
  NOR2_X1 U157 ( .A1(S[1]), .A2(S[2]), .ZN(n309) );
  INV_X1 U158 ( .A(S[2]), .ZN(n312) );
  NAND4_X2 U159 ( .A1(n316), .A2(n315), .A3(n314), .A4(n313), .ZN(Y[0]) );
  INV_X1 U160 ( .A(D[1]), .ZN(n317) );
  INV_X1 U161 ( .A(B[1]), .ZN(n318) );
  NOR2_X1 U162 ( .A1(n320), .A2(n319), .ZN(n323) );
  NAND2_X1 U163 ( .A1(A[1]), .A2(n396), .ZN(n322) );
  AOI22_X1 U164 ( .A1(C[1]), .A2(n247), .B1(E[1]), .B2(n245), .ZN(n321) );
  NAND3_X1 U165 ( .A1(n323), .A2(n322), .A3(n321), .ZN(Y[1]) );
  INV_X1 U166 ( .A(D[2]), .ZN(n324) );
  INV_X1 U167 ( .A(B[2]), .ZN(n325) );
  NOR2_X1 U168 ( .A1(n327), .A2(n326), .ZN(n330) );
  NAND2_X1 U169 ( .A1(A[2]), .A2(n396), .ZN(n329) );
  AOI22_X1 U170 ( .A1(C[2]), .A2(n248), .B1(E[2]), .B2(n245), .ZN(n328) );
  NAND3_X1 U171 ( .A1(n330), .A2(n329), .A3(n328), .ZN(Y[2]) );
  INV_X1 U172 ( .A(D[3]), .ZN(n331) );
  INV_X1 U173 ( .A(B[3]), .ZN(n332) );
  NOR2_X1 U174 ( .A1(n334), .A2(n333), .ZN(n337) );
  NAND2_X1 U175 ( .A1(A[3]), .A2(n239), .ZN(n336) );
  AOI22_X1 U176 ( .A1(C[3]), .A2(n248), .B1(E[3]), .B2(n245), .ZN(n335) );
  NAND3_X1 U177 ( .A1(n337), .A2(n336), .A3(n335), .ZN(Y[3]) );
  INV_X1 U178 ( .A(D[4]), .ZN(n338) );
  NOR2_X1 U179 ( .A1(n340), .A2(n339), .ZN(n343) );
  NAND2_X1 U180 ( .A1(A[4]), .A2(n239), .ZN(n342) );
  AOI22_X1 U181 ( .A1(C[4]), .A2(n247), .B1(E[4]), .B2(n245), .ZN(n341) );
  NOR2_X1 U182 ( .A1(n345), .A2(n344), .ZN(n348) );
  NAND2_X1 U183 ( .A1(A[5]), .A2(n239), .ZN(n347) );
  AOI22_X1 U184 ( .A1(C[5]), .A2(n247), .B1(E[5]), .B2(n245), .ZN(n346) );
  NAND3_X1 U185 ( .A1(n348), .A2(n347), .A3(n346), .ZN(Y[5]) );
  NOR2_X1 U186 ( .A1(n350), .A2(n349), .ZN(n353) );
  NAND2_X1 U187 ( .A1(A[6]), .A2(n396), .ZN(n352) );
  AOI22_X1 U188 ( .A1(C[6]), .A2(n247), .B1(E[6]), .B2(n245), .ZN(n351) );
  NAND3_X1 U189 ( .A1(n353), .A2(n352), .A3(n351), .ZN(Y[6]) );
  NOR2_X1 U190 ( .A1(n355), .A2(n354), .ZN(n358) );
  NAND2_X1 U191 ( .A1(A[7]), .A2(n239), .ZN(n357) );
  AOI22_X1 U192 ( .A1(C[7]), .A2(n247), .B1(E[7]), .B2(n245), .ZN(n356) );
  NAND3_X1 U193 ( .A1(n358), .A2(n357), .A3(n356), .ZN(Y[7]) );
  NOR2_X1 U194 ( .A1(n360), .A2(n359), .ZN(n363) );
  NAND2_X1 U195 ( .A1(A[8]), .A2(n239), .ZN(n362) );
  AOI22_X1 U196 ( .A1(C[8]), .A2(n247), .B1(E[8]), .B2(n245), .ZN(n361) );
  NAND3_X1 U197 ( .A1(n363), .A2(n362), .A3(n361), .ZN(Y[8]) );
  NOR2_X1 U198 ( .A1(n365), .A2(n364), .ZN(n368) );
  NAND2_X1 U199 ( .A1(A[9]), .A2(n239), .ZN(n367) );
  AOI22_X1 U200 ( .A1(C[9]), .A2(n247), .B1(E[9]), .B2(n245), .ZN(n366) );
  NAND3_X1 U201 ( .A1(n368), .A2(n367), .A3(n366), .ZN(Y[9]) );
  NOR2_X1 U202 ( .A1(n370), .A2(n369), .ZN(n373) );
  NAND2_X1 U203 ( .A1(A[10]), .A2(n396), .ZN(n372) );
  AOI22_X1 U204 ( .A1(C[10]), .A2(n247), .B1(E[10]), .B2(n245), .ZN(n371) );
  NAND3_X1 U205 ( .A1(n373), .A2(n372), .A3(n371), .ZN(Y[10]) );
  NOR2_X1 U206 ( .A1(n375), .A2(n374), .ZN(n378) );
  NAND2_X1 U207 ( .A1(A[11]), .A2(n239), .ZN(n377) );
  AOI22_X1 U208 ( .A1(C[11]), .A2(n247), .B1(E[11]), .B2(n245), .ZN(n376) );
  NAND3_X1 U209 ( .A1(n378), .A2(n377), .A3(n376), .ZN(Y[11]) );
  NOR2_X1 U210 ( .A1(n380), .A2(n379), .ZN(n383) );
  NAND2_X1 U211 ( .A1(A[12]), .A2(n239), .ZN(n382) );
  AOI22_X1 U212 ( .A1(C[12]), .A2(n247), .B1(E[12]), .B2(n245), .ZN(n381) );
  NAND3_X1 U213 ( .A1(n383), .A2(n382), .A3(n381), .ZN(Y[12]) );
  NOR2_X1 U214 ( .A1(n385), .A2(n384), .ZN(n388) );
  NAND2_X1 U215 ( .A1(A[13]), .A2(n239), .ZN(n387) );
  AOI22_X1 U216 ( .A1(C[13]), .A2(n247), .B1(E[13]), .B2(n245), .ZN(n386) );
  NAND3_X1 U217 ( .A1(n388), .A2(n387), .A3(n386), .ZN(Y[13]) );
  NOR2_X1 U218 ( .A1(n390), .A2(n389), .ZN(n393) );
  NAND2_X1 U219 ( .A1(A[14]), .A2(n239), .ZN(n392) );
  AOI22_X1 U220 ( .A1(C[14]), .A2(n247), .B1(E[14]), .B2(n245), .ZN(n391) );
  NAND3_X1 U221 ( .A1(n393), .A2(n392), .A3(n391), .ZN(Y[14]) );
  NOR2_X1 U222 ( .A1(n395), .A2(n394), .ZN(n399) );
  NAND2_X1 U223 ( .A1(A[15]), .A2(n239), .ZN(n398) );
  AOI22_X1 U224 ( .A1(C[15]), .A2(n247), .B1(E[15]), .B2(n245), .ZN(n397) );
  NAND3_X1 U225 ( .A1(n399), .A2(n398), .A3(n397), .ZN(Y[15]) );
  NAND2_X1 U226 ( .A1(E[16]), .A2(n245), .ZN(n405) );
  INV_X1 U227 ( .A(A[16]), .ZN(n400) );
  OAI22_X1 U228 ( .A1(n252), .A2(n303), .B1(n250), .B2(n300), .ZN(n401) );
  NOR2_X1 U229 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND3_X1 U230 ( .A1(n405), .A2(n404), .A3(n403), .ZN(Y[16]) );
  NAND2_X1 U231 ( .A1(C[17]), .A2(n248), .ZN(n410) );
  INV_X1 U232 ( .A(A[17]), .ZN(n406) );
  OAI22_X1 U233 ( .A1(n252), .A2(n305), .B1(n250), .B2(n302), .ZN(n407) );
  NOR2_X1 U234 ( .A1(n408), .A2(n407), .ZN(n409) );
  NAND3_X1 U235 ( .A1(n411), .A2(n410), .A3(n409), .ZN(Y[17]) );
  NAND2_X1 U236 ( .A1(E[18]), .A2(n245), .ZN(n417) );
  INV_X1 U237 ( .A(A[18]), .ZN(n412) );
  OAI22_X1 U238 ( .A1(n252), .A2(n307), .B1(n250), .B2(n304), .ZN(n413) );
  NOR2_X1 U239 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND3_X1 U240 ( .A1(n417), .A2(n416), .A3(n415), .ZN(Y[18]) );
  INV_X1 U241 ( .A(A[19]), .ZN(n418) );
  OAI22_X1 U242 ( .A1(n252), .A2(n269), .B1(n250), .B2(n306), .ZN(n419) );
  NOR2_X1 U243 ( .A1(n420), .A2(n419), .ZN(n421) );
  NAND3_X1 U244 ( .A1(n423), .A2(n422), .A3(n421), .ZN(Y[19]) );
  INV_X1 U245 ( .A(A[20]), .ZN(n424) );
  OAI22_X1 U246 ( .A1(n252), .A2(n270), .B1(n250), .B2(n257), .ZN(n425) );
  NOR2_X1 U247 ( .A1(n426), .A2(n425), .ZN(n427) );
  INV_X1 U248 ( .A(A[21]), .ZN(n430) );
  OAI22_X1 U249 ( .A1(n252), .A2(n271), .B1(n250), .B2(n258), .ZN(n431) );
  NOR2_X1 U250 ( .A1(n432), .A2(n431), .ZN(n433) );
  NAND3_X1 U251 ( .A1(n435), .A2(n434), .A3(n433), .ZN(Y[21]) );
  INV_X1 U252 ( .A(A[22]), .ZN(n436) );
  OAI22_X1 U253 ( .A1(n252), .A2(n272), .B1(n250), .B2(n259), .ZN(n437) );
  NOR2_X1 U254 ( .A1(n438), .A2(n437), .ZN(n439) );
  NAND3_X1 U255 ( .A1(n441), .A2(n440), .A3(n439), .ZN(Y[22]) );
  INV_X1 U256 ( .A(A[23]), .ZN(n442) );
  OAI22_X1 U257 ( .A1(n252), .A2(n273), .B1(n250), .B2(n260), .ZN(n443) );
  NOR2_X1 U258 ( .A1(n444), .A2(n443), .ZN(n445) );
  NAND3_X1 U259 ( .A1(n447), .A2(n446), .A3(n445), .ZN(Y[23]) );
  INV_X1 U260 ( .A(A[24]), .ZN(n448) );
  OAI22_X1 U261 ( .A1(n252), .A2(n274), .B1(n250), .B2(n261), .ZN(n449) );
  NOR2_X1 U262 ( .A1(n450), .A2(n449), .ZN(n451) );
  NAND3_X1 U263 ( .A1(n453), .A2(n452), .A3(n451), .ZN(Y[24]) );
  INV_X1 U264 ( .A(A[25]), .ZN(n454) );
  OAI22_X1 U265 ( .A1(n252), .A2(n275), .B1(n250), .B2(n262), .ZN(n455) );
  NOR2_X1 U266 ( .A1(n456), .A2(n455), .ZN(n457) );
  NAND3_X1 U267 ( .A1(n459), .A2(n458), .A3(n457), .ZN(Y[25]) );
  INV_X1 U268 ( .A(A[26]), .ZN(n460) );
  OAI22_X1 U269 ( .A1(n252), .A2(n276), .B1(n250), .B2(n263), .ZN(n461) );
  NOR2_X1 U270 ( .A1(n462), .A2(n461), .ZN(n463) );
  NAND3_X1 U271 ( .A1(n465), .A2(n464), .A3(n463), .ZN(Y[26]) );
  INV_X1 U272 ( .A(A[27]), .ZN(n466) );
  OAI22_X1 U273 ( .A1(n252), .A2(n277), .B1(n250), .B2(n264), .ZN(n467) );
  NOR2_X1 U274 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND3_X1 U275 ( .A1(n471), .A2(n470), .A3(n469), .ZN(Y[27]) );
  INV_X1 U276 ( .A(A[28]), .ZN(n472) );
  OAI22_X1 U277 ( .A1(n252), .A2(n278), .B1(n250), .B2(n265), .ZN(n473) );
  NOR2_X1 U278 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND3_X1 U279 ( .A1(n477), .A2(n476), .A3(n475), .ZN(Y[28]) );
  INV_X1 U280 ( .A(A[29]), .ZN(n478) );
  OAI22_X1 U281 ( .A1(n252), .A2(n279), .B1(n250), .B2(n266), .ZN(n479) );
  NOR2_X1 U282 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND3_X1 U283 ( .A1(n483), .A2(n482), .A3(n481), .ZN(Y[29]) );
  INV_X1 U284 ( .A(A[30]), .ZN(n484) );
  OAI22_X1 U285 ( .A1(n252), .A2(n280), .B1(n250), .B2(n267), .ZN(n485) );
  NOR2_X1 U286 ( .A1(n486), .A2(n485), .ZN(n487) );
  NAND3_X1 U287 ( .A1(n489), .A2(n488), .A3(n487), .ZN(Y[30]) );
  INV_X1 U288 ( .A(A[31]), .ZN(n490) );
  OAI22_X1 U289 ( .A1(n252), .A2(n281), .B1(n250), .B2(n268), .ZN(n492) );
  NOR2_X1 U290 ( .A1(n493), .A2(n492), .ZN(n494) );
  NAND3_X1 U291 ( .A1(n496), .A2(n495), .A3(n494), .ZN(Y[31]) );
endmodule


module Boothencoder_6 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   n8, n10, n11, n12;

  BUF_X1 U1 ( .A(n12), .Z(n8) );
  OAI21_X1 U2 ( .B1(B[0]), .B2(B[1]), .A(n12), .ZN(n11) );
  NAND2_X1 U3 ( .A1(B[1]), .A2(B[0]), .ZN(n12) );
  AND3_X1 U4 ( .A1(n11), .A2(B[2]), .A3(n8), .ZN(S[2]) );
  AOI21_X1 U5 ( .B1(n8), .B2(n11), .A(B[2]), .ZN(S[0]) );
  MUX2_X1 U6 ( .A(n8), .B(n11), .S(B[2]), .Z(n10) );
  INV_X1 U7 ( .A(n10), .ZN(S[1]) );
endmodule


module p4adder_N32_7 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;
  wire   n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;
  wire   [8:0] C;
  assign n1 = A[11];
  assign n4 = A[15];
  assign n5 = B[3];
  assign n6 = A[1];
  assign n7 = A[0];
  assign n8 = A[3];
  assign n9 = A[5];
  assign n10 = B[5];
  assign n11 = B[6];
  assign n12 = A[10];
  assign n13 = A[6];
  assign n14 = B[11];
  assign n15 = B[14];
  assign n16 = B[7];
  assign n17 = A[7];

  CarryGen_N32_7 Cgen ( .A({A[31:16], n4, A[14:12], n1, n12, A[9:8], n17, n13, 
        n9, A[4], n8, A[2], n6, n37}), .B({B[31:21], n18, B[19:15], n15, 
        B[13:12], n14, B[10:8], n16, n11, n10, n22, n5, B[2:1], n23}), .Cin(
        Cin), .C(C) );
  SumGen_N32_7 Sgen ( .A({A[31:16], n39, A[14:12], n40, n12, A[9:8], n38, n29, 
        n28, A[4], n35, n20, n25, n21}), .B({B[31:21], n18, B[19:16], n27, n32, 
        B[13:12], n33, B[10:8], n36, n30, n34, n26, n41, n19, n24, n31}), .C(C), .S(S), .Cout(Cout) );
  BUF_X2 U1 ( .A(B[20]), .Z(n18) );
  CLKBUF_X1 U2 ( .A(n16), .Z(n36) );
  CLKBUF_X1 U3 ( .A(n5), .Z(n41) );
  CLKBUF_X1 U4 ( .A(n17), .Z(n38) );
  BUF_X2 U5 ( .A(B[2]), .Z(n19) );
  BUF_X1 U6 ( .A(A[2]), .Z(n20) );
  CLKBUF_X3 U7 ( .A(n7), .Z(n21) );
  CLKBUF_X1 U8 ( .A(n7), .Z(n37) );
  CLKBUF_X1 U9 ( .A(B[4]), .Z(n22) );
  BUF_X2 U10 ( .A(B[4]), .Z(n26) );
  CLKBUF_X1 U11 ( .A(B[0]), .Z(n23) );
  BUF_X2 U12 ( .A(B[1]), .Z(n24) );
  BUF_X2 U13 ( .A(n6), .Z(n25) );
  CLKBUF_X1 U14 ( .A(B[15]), .Z(n27) );
  BUF_X2 U15 ( .A(n9), .Z(n28) );
  BUF_X1 U16 ( .A(n13), .Z(n29) );
  BUF_X1 U17 ( .A(n11), .Z(n30) );
  BUF_X2 U18 ( .A(B[0]), .Z(n31) );
  BUF_X1 U19 ( .A(n15), .Z(n32) );
  CLKBUF_X1 U20 ( .A(n14), .Z(n33) );
  BUF_X2 U21 ( .A(n10), .Z(n34) );
  CLKBUF_X1 U22 ( .A(n8), .Z(n35) );
  CLKBUF_X1 U23 ( .A(n4), .Z(n39) );
  CLKBUF_X1 U24 ( .A(n1), .Z(n40) );
endmodule


module mux51_generic_N32_7 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   net227453, net227454, net227465, net227476, net227484, net227488,
         net227489, net227494, net227502, net227514, net227530, net227532,
         net227551, net227557, net227604, net227607, net227609, net227610,
         net227611, net227624, net227626, net227627, net227636, net227640,
         net227644, net227647, net227648, net232336, net232999, net239666,
         net239669, net239670, net239684, net239854, net239905, net240023,
         net233271, net241293, net241372, net241371, net241471, net239677,
         net233026, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446;

  AND2_X1 U2 ( .A1(n300), .A2(net239854), .ZN(n345) );
  AND2_X1 U3 ( .A1(S[0]), .A2(D[3]), .ZN(n300) );
  INV_X1 U4 ( .A(n314), .ZN(n301) );
  OR2_X2 U5 ( .A1(n312), .A2(net227636), .ZN(n314) );
  AND2_X2 U6 ( .A1(n313), .A2(n308), .ZN(net239670) );
  AOI211_X4 U7 ( .C1(E[16]), .C2(net232336), .A(n396), .B(n395), .ZN(n397) );
  NAND4_X1 U8 ( .A1(net227624), .A2(n342), .A3(net227626), .A4(net227627), 
        .ZN(Y[2]) );
  BUF_X1 U9 ( .A(net239666), .Z(n311) );
  INV_X2 U10 ( .A(net227454), .ZN(net227465) );
  INV_X2 U11 ( .A(net241371), .ZN(net227488) );
  INV_X1 U12 ( .A(net227636), .ZN(n302) );
  INV_X1 U13 ( .A(net239854), .ZN(n303) );
  AND2_X1 U14 ( .A1(net227607), .A2(n327), .ZN(n304) );
  BUF_X2 U15 ( .A(net239669), .Z(net232336) );
  AND3_X1 U16 ( .A1(n381), .A2(n379), .A3(n380), .ZN(n305) );
  AND3_X1 U17 ( .A1(n382), .A2(n383), .A3(n384), .ZN(n306) );
  NAND2_X1 U18 ( .A1(n385), .A2(n306), .ZN(Y[13]) );
  INV_X1 U19 ( .A(n325), .ZN(n307) );
  AND2_X2 U20 ( .A1(n312), .A2(net241293), .ZN(n330) );
  NAND4_X1 U21 ( .A1(n363), .A2(n364), .A3(n365), .A4(n362), .ZN(Y[8]) );
  BUF_X1 U22 ( .A(net239677), .Z(n309) );
  BUF_X1 U23 ( .A(net239677), .Z(n308) );
  BUF_X1 U24 ( .A(net239677), .Z(net241293) );
  AND2_X1 U25 ( .A1(E[6]), .A2(net239669), .ZN(n310) );
  NOR2_X1 U26 ( .A1(n310), .A2(n353), .ZN(n357) );
  AOI22_X1 U27 ( .A1(E[1]), .A2(n304), .B1(n322), .B2(B[1]), .ZN(n316) );
  AND2_X2 U28 ( .A1(net227607), .A2(n327), .ZN(net239669) );
  AND2_X1 U29 ( .A1(n325), .A2(n308), .ZN(net239684) );
  AND2_X1 U30 ( .A1(n325), .A2(net241293), .ZN(net232999) );
  INV_X1 U31 ( .A(n321), .ZN(n313) );
  INV_X1 U32 ( .A(n321), .ZN(n312) );
  OR2_X1 U33 ( .A1(net233271), .A2(net227636), .ZN(net227453) );
  NAND4_X1 U34 ( .A1(n316), .A2(n318), .A3(n317), .A4(n319), .ZN(Y[1]) );
  NAND2_X1 U35 ( .A1(C[1]), .A2(net233026), .ZN(n319) );
  NAND2_X1 U36 ( .A1(A[1]), .A2(n320), .ZN(n317) );
  NAND2_X1 U37 ( .A1(net239905), .A2(D[1]), .ZN(n318) );
  AND2_X1 U38 ( .A1(n312), .A2(n309), .ZN(net233026) );
  NAND2_X1 U39 ( .A1(net233026), .A2(C[2]), .ZN(net227627) );
  NOR2_X1 U40 ( .A1(S[0]), .A2(S[2]), .ZN(net239677) );
  INV_X1 U41 ( .A(S[1]), .ZN(n321) );
  INV_X1 U42 ( .A(n321), .ZN(net233271) );
  AND2_X1 U43 ( .A1(net241293), .A2(n325), .ZN(n320) );
  AND2_X1 U44 ( .A1(n320), .A2(A[14]), .ZN(net227557) );
  AOI22_X1 U45 ( .A1(E[4]), .A2(net239669), .B1(A[4]), .B2(n320), .ZN(
        net227609) );
  INV_X1 U46 ( .A(n324), .ZN(n325) );
  BUF_X1 U47 ( .A(S[1]), .Z(n324) );
  INV_X1 U48 ( .A(n324), .ZN(net227607) );
  AND2_X1 U49 ( .A1(n315), .A2(n313), .ZN(n323) );
  NAND2_X1 U50 ( .A1(net239905), .A2(D[2]), .ZN(net227626) );
  INV_X1 U51 ( .A(net227636), .ZN(n315) );
  AND2_X1 U52 ( .A1(n315), .A2(n312), .ZN(net241471) );
  AND2_X1 U53 ( .A1(n302), .A2(n313), .ZN(net239905) );
  NOR2_X1 U54 ( .A1(net233271), .A2(net227636), .ZN(n322) );
  AOI22_X1 U55 ( .A1(E[2]), .A2(net239666), .B1(n322), .B2(B[2]), .ZN(
        net227624) );
  NAND3_X1 U56 ( .A1(net227604), .A2(n351), .A3(n352), .ZN(Y[5]) );
  INV_X1 U57 ( .A(n323), .ZN(net241372) );
  INV_X1 U58 ( .A(net241471), .ZN(net241371) );
  NAND3_X1 U59 ( .A1(n355), .A2(n356), .A3(n357), .ZN(Y[6]) );
  NAND2_X1 U60 ( .A1(n323), .A2(D[4]), .ZN(net227611) );
  AOI22_X1 U61 ( .A1(D[5]), .A2(net241471), .B1(C[5]), .B2(n330), .ZN(
        net227604) );
  NAND3_X1 U62 ( .A1(net227647), .A2(net227648), .A3(net233271), .ZN(net227644) );
  NAND2_X1 U63 ( .A1(net227551), .A2(B[4]), .ZN(net227610) );
  NAND3_X2 U64 ( .A1(n404), .A2(n403), .A3(n402), .ZN(Y[17]) );
  NAND2_X2 U65 ( .A1(n378), .A2(n305), .ZN(Y[12]) );
  NAND4_X2 U66 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .ZN(Y[10]) );
  NAND3_X2 U67 ( .A1(n389), .A2(n390), .A3(n391), .ZN(Y[14]) );
  NAND4_X2 U68 ( .A1(n369), .A2(n366), .A3(n367), .A4(n368), .ZN(Y[9]) );
  INV_X1 U69 ( .A(S[2]), .ZN(net240023) );
  AND2_X1 U70 ( .A1(D[6]), .A2(n323), .ZN(n326) );
  NOR2_X1 U71 ( .A1(n326), .A2(n354), .ZN(n355) );
  NAND2_X1 U72 ( .A1(n349), .A2(n348), .ZN(Y[3]) );
  INV_X1 U73 ( .A(S[2]), .ZN(net239854) );
  AND2_X1 U74 ( .A1(C[6]), .A2(n330), .ZN(n354) );
  AND2_X1 U75 ( .A1(net227607), .A2(n327), .ZN(net239666) );
  AND2_X1 U76 ( .A1(net227640), .A2(S[2]), .ZN(n327) );
  AOI22_X1 U77 ( .A1(A[28]), .A2(net227465), .B1(B[28]), .B2(net227502), .ZN(
        n437) );
  NAND2_X1 U78 ( .A1(E[28]), .A2(n311), .ZN(n436) );
  AOI22_X1 U79 ( .A1(A[29]), .A2(net227465), .B1(B[29]), .B2(net227502), .ZN(
        n440) );
  NAND2_X1 U80 ( .A1(E[29]), .A2(net232336), .ZN(n439) );
  AOI22_X1 U81 ( .A1(A[22]), .A2(net227465), .B1(B[22]), .B2(net227502), .ZN(
        n419) );
  AOI22_X1 U82 ( .A1(A[23]), .A2(net227465), .B1(B[23]), .B2(net227502), .ZN(
        n422) );
  NAND2_X1 U83 ( .A1(E[23]), .A2(net232336), .ZN(n421) );
  AOI22_X1 U84 ( .A1(A[25]), .A2(net227489), .B1(B[25]), .B2(net227532), .ZN(
        n428) );
  NAND2_X1 U85 ( .A1(E[25]), .A2(net232336), .ZN(n427) );
  AOI22_X1 U86 ( .A1(A[27]), .A2(net227465), .B1(B[27]), .B2(net227532), .ZN(
        n434) );
  NAND2_X1 U87 ( .A1(E[27]), .A2(net232336), .ZN(n433) );
  AOI22_X1 U88 ( .A1(A[18]), .A2(net227465), .B1(B[18]), .B2(net227532), .ZN(
        n407) );
  AOI22_X1 U89 ( .A1(D[18]), .A2(net227488), .B1(C[18]), .B2(n328), .ZN(n405)
         );
  AOI22_X1 U90 ( .A1(A[24]), .A2(net227465), .B1(B[24]), .B2(net227502), .ZN(
        n425) );
  NAND2_X1 U91 ( .A1(E[24]), .A2(net232336), .ZN(n424) );
  AOI22_X1 U92 ( .A1(D[24]), .A2(net227494), .B1(C[24]), .B2(net239670), .ZN(
        n423) );
  AOI22_X1 U93 ( .A1(A[21]), .A2(net227465), .B1(B[21]), .B2(net227502), .ZN(
        n416) );
  NAND2_X1 U94 ( .A1(E[21]), .A2(n311), .ZN(n415) );
  AOI22_X1 U95 ( .A1(D[21]), .A2(net227476), .B1(C[21]), .B2(n330), .ZN(n414)
         );
  AOI22_X1 U96 ( .A1(A[26]), .A2(net227489), .B1(B[26]), .B2(net227502), .ZN(
        n431) );
  NAND2_X1 U97 ( .A1(E[26]), .A2(net232336), .ZN(n430) );
  AOI22_X1 U98 ( .A1(D[26]), .A2(net227488), .B1(C[26]), .B2(n330), .ZN(n429)
         );
  AOI22_X1 U99 ( .A1(A[19]), .A2(net227489), .B1(B[19]), .B2(net227502), .ZN(
        n410) );
  AOI22_X1 U100 ( .A1(D[19]), .A2(net227488), .B1(C[19]), .B2(n330), .ZN(n408)
         );
  AOI22_X1 U101 ( .A1(A[20]), .A2(net227489), .B1(B[20]), .B2(net227502), .ZN(
        n413) );
  AOI22_X1 U102 ( .A1(D[20]), .A2(net227488), .B1(C[20]), .B2(n329), .ZN(n411)
         );
  AND2_X1 U103 ( .A1(net239684), .A2(A[16]), .ZN(n396) );
  AND2_X1 U104 ( .A1(net232999), .A2(A[17]), .ZN(n401) );
  AOI22_X1 U105 ( .A1(A[31]), .A2(net227465), .B1(B[31]), .B2(net227532), .ZN(
        n446) );
  AOI22_X1 U106 ( .A1(A[30]), .A2(net227489), .B1(B[30]), .B2(net227532), .ZN(
        n443) );
  NAND2_X1 U107 ( .A1(E[30]), .A2(net232336), .ZN(n442) );
  AOI22_X1 U108 ( .A1(D[30]), .A2(net227488), .B1(C[30]), .B2(net239670), .ZN(
        n441) );
  NOR2_X1 U109 ( .A1(n340), .A2(n341), .ZN(Y[0]) );
  NAND4_X1 U110 ( .A1(n361), .A2(n359), .A3(n360), .A4(n358), .ZN(Y[7]) );
  NAND3_X1 U111 ( .A1(n394), .A2(n393), .A3(n392), .ZN(Y[15]) );
  AND2_X1 U112 ( .A1(n312), .A2(n309), .ZN(n329) );
  AND2_X1 U113 ( .A1(n308), .A2(n313), .ZN(n328) );
  AOI21_X1 U114 ( .B1(A[3]), .B2(n308), .A(n344), .ZN(n347) );
  AOI211_X1 U115 ( .C1(E[17]), .C2(n311), .A(n401), .B(n400), .ZN(n402) );
  AOI22_X1 U116 ( .A1(D[31]), .A2(net227488), .B1(C[31]), .B2(n328), .ZN(n444)
         );
  AOI22_X1 U117 ( .A1(D[29]), .A2(net227530), .B1(C[29]), .B2(n328), .ZN(n438)
         );
  AOI22_X1 U118 ( .A1(D[28]), .A2(net227488), .B1(C[28]), .B2(n329), .ZN(n435)
         );
  AOI22_X1 U119 ( .A1(D[27]), .A2(net227488), .B1(C[27]), .B2(n328), .ZN(n432)
         );
  AOI22_X1 U120 ( .A1(D[25]), .A2(net227488), .B1(C[25]), .B2(n328), .ZN(n426)
         );
  AOI22_X1 U121 ( .A1(D[23]), .A2(net227488), .B1(C[23]), .B2(n329), .ZN(n420)
         );
  AOI22_X1 U122 ( .A1(D[22]), .A2(net227476), .B1(C[22]), .B2(n328), .ZN(n417)
         );
  NAND2_X1 U123 ( .A1(C[14]), .A2(n330), .ZN(n390) );
  NAND4_X2 U124 ( .A1(net227609), .A2(net227610), .A3(net227611), .A4(n350), 
        .ZN(Y[4]) );
  NAND2_X1 U125 ( .A1(C[17]), .A2(net239670), .ZN(n403) );
  INV_X1 U126 ( .A(net232999), .ZN(net227454) );
  INV_X1 U127 ( .A(net241371), .ZN(net227476) );
  INV_X1 U128 ( .A(net241372), .ZN(net227530) );
  AOI21_X1 U129 ( .B1(C[3]), .B2(n309), .A(n345), .ZN(n346) );
  NAND2_X1 U130 ( .A1(C[16]), .A2(n329), .ZN(n398) );
  NAND2_X1 U131 ( .A1(E[31]), .A2(n311), .ZN(n445) );
  NAND2_X1 U132 ( .A1(E[22]), .A2(net232336), .ZN(n418) );
  NAND2_X1 U133 ( .A1(E[20]), .A2(net232336), .ZN(n412) );
  NAND2_X1 U134 ( .A1(E[18]), .A2(net232336), .ZN(n406) );
  NAND2_X1 U135 ( .A1(E[19]), .A2(net232336), .ZN(n409) );
  AOI22_X1 U136 ( .A1(B[15]), .A2(net227514), .B1(E[15]), .B2(net232336), .ZN(
        n392) );
  INV_X1 U137 ( .A(net241372), .ZN(net227494) );
  INV_X1 U138 ( .A(net227453), .ZN(net227484) );
  INV_X1 U139 ( .A(n314), .ZN(net227502) );
  INV_X1 U140 ( .A(n314), .ZN(net227514) );
  INV_X1 U141 ( .A(n314), .ZN(net227532) );
  NOR2_X1 U142 ( .A1(n314), .A2(n331), .ZN(n400) );
  NOR2_X1 U143 ( .A1(n314), .A2(n333), .ZN(n395) );
  INV_X1 U144 ( .A(net227453), .ZN(net227551) );
  NOR2_X1 U145 ( .A1(n314), .A2(n332), .ZN(n353) );
  AOI22_X1 U146 ( .A1(D[15]), .A2(net227488), .B1(C[15]), .B2(n328), .ZN(n394)
         );
  NAND2_X1 U147 ( .A1(A[15]), .A2(net227489), .ZN(n393) );
  NAND2_X1 U148 ( .A1(A[5]), .A2(net239684), .ZN(n351) );
  AOI22_X1 U149 ( .A1(B[5]), .A2(net227484), .B1(net239669), .B2(E[5]), .ZN(
        n352) );
  NAND2_X1 U150 ( .A1(S[0]), .A2(net240023), .ZN(net227636) );
  INV_X1 U151 ( .A(net227454), .ZN(net227489) );
  INV_X1 U152 ( .A(B[17]), .ZN(n331) );
  INV_X1 U153 ( .A(B[6]), .ZN(n332) );
  INV_X1 U154 ( .A(B[16]), .ZN(n333) );
  INV_X1 U155 ( .A(B[0]), .ZN(n334) );
  OAI21_X1 U156 ( .B1(n334), .B2(n303), .A(S[0]), .ZN(n335) );
  AOI21_X1 U157 ( .B1(n307), .B2(net239854), .A(n335), .ZN(n341) );
  INV_X1 U158 ( .A(A[0]), .ZN(n336) );
  INV_X1 U159 ( .A(S[0]), .ZN(net227640) );
  NAND2_X1 U160 ( .A1(n336), .A2(n309), .ZN(n339) );
  NAND2_X1 U161 ( .A1(S[0]), .A2(D[0]), .ZN(net227647) );
  NAND3_X1 U162 ( .A1(net227640), .A2(net239854), .A3(C[0]), .ZN(net227648) );
  INV_X1 U163 ( .A(E[0]), .ZN(n337) );
  NAND2_X1 U164 ( .A1(n303), .A2(n337), .ZN(n338) );
  OAI211_X1 U165 ( .C1(n339), .C2(n313), .A(net227644), .B(n338), .ZN(n340) );
  NAND2_X1 U166 ( .A1(A[2]), .A2(net232999), .ZN(n342) );
  NAND2_X1 U167 ( .A1(net227484), .A2(B[3]), .ZN(n349) );
  NAND2_X1 U168 ( .A1(S[2]), .A2(E[3]), .ZN(n343) );
  NOR2_X1 U169 ( .A1(n343), .A2(S[0]), .ZN(n344) );
  MUX2_X1 U170 ( .A(n347), .B(n346), .S(n307), .Z(n348) );
  NAND2_X1 U171 ( .A1(C[4]), .A2(net239670), .ZN(n350) );
  NAND2_X1 U172 ( .A1(A[6]), .A2(net239684), .ZN(n356) );
  AOI22_X1 U173 ( .A1(E[7]), .A2(net239669), .B1(net227551), .B2(B[7]), .ZN(
        n361) );
  NAND2_X1 U174 ( .A1(A[7]), .A2(net239684), .ZN(n360) );
  NAND2_X1 U175 ( .A1(D[7]), .A2(net241471), .ZN(n359) );
  NAND2_X1 U176 ( .A1(C[7]), .A2(n329), .ZN(n358) );
  AOI22_X1 U177 ( .A1(E[8]), .A2(n311), .B1(n301), .B2(B[8]), .ZN(n365) );
  NAND2_X1 U178 ( .A1(A[8]), .A2(net239684), .ZN(n364) );
  NAND2_X1 U179 ( .A1(D[8]), .A2(net227530), .ZN(n363) );
  NAND2_X1 U180 ( .A1(C[8]), .A2(net239670), .ZN(n362) );
  AOI22_X1 U181 ( .A1(E[9]), .A2(n311), .B1(B[9]), .B2(net227514), .ZN(n369)
         );
  NAND2_X1 U182 ( .A1(A[9]), .A2(net239684), .ZN(n368) );
  NAND2_X1 U183 ( .A1(D[9]), .A2(net227494), .ZN(n367) );
  NAND2_X1 U184 ( .A1(C[9]), .A2(n328), .ZN(n366) );
  AOI22_X1 U185 ( .A1(E[10]), .A2(net232336), .B1(B[10]), .B2(net227532), .ZN(
        n373) );
  NAND2_X1 U186 ( .A1(A[10]), .A2(net232999), .ZN(n372) );
  NAND2_X1 U187 ( .A1(D[10]), .A2(net227476), .ZN(n371) );
  NAND2_X1 U188 ( .A1(C[10]), .A2(n329), .ZN(n370) );
  AOI22_X1 U189 ( .A1(E[11]), .A2(net232336), .B1(B[11]), .B2(net227514), .ZN(
        n377) );
  NAND2_X1 U190 ( .A1(A[11]), .A2(net232999), .ZN(n376) );
  NAND2_X1 U191 ( .A1(D[11]), .A2(net227494), .ZN(n375) );
  NAND2_X1 U192 ( .A1(C[11]), .A2(n330), .ZN(n374) );
  NAND4_X1 U193 ( .A1(n377), .A2(n376), .A3(n375), .A4(n374), .ZN(Y[11]) );
  AOI22_X1 U194 ( .A1(E[12]), .A2(net232336), .B1(net227502), .B2(B[12]), .ZN(
        n381) );
  NAND2_X1 U195 ( .A1(A[12]), .A2(net232999), .ZN(n380) );
  NAND2_X1 U196 ( .A1(D[12]), .A2(net227530), .ZN(n379) );
  NAND2_X1 U197 ( .A1(C[12]), .A2(n328), .ZN(n378) );
  AOI22_X1 U198 ( .A1(E[13]), .A2(net232336), .B1(B[13]), .B2(net227532), .ZN(
        n385) );
  NAND2_X1 U199 ( .A1(A[13]), .A2(net239684), .ZN(n384) );
  NAND2_X1 U200 ( .A1(D[13]), .A2(net227476), .ZN(n383) );
  NAND2_X1 U201 ( .A1(C[13]), .A2(net239670), .ZN(n382) );
  NAND2_X1 U202 ( .A1(D[14]), .A2(net227488), .ZN(n391) );
  NAND2_X1 U203 ( .A1(B[14]), .A2(net227514), .ZN(n387) );
  NAND2_X1 U204 ( .A1(E[14]), .A2(n311), .ZN(n386) );
  NAND2_X1 U205 ( .A1(n386), .A2(n387), .ZN(n388) );
  NOR2_X1 U206 ( .A1(net227557), .A2(n388), .ZN(n389) );
  NAND2_X1 U207 ( .A1(D[16]), .A2(net227488), .ZN(n399) );
  NAND3_X1 U208 ( .A1(n399), .A2(n398), .A3(n397), .ZN(Y[16]) );
  NAND2_X1 U209 ( .A1(D[17]), .A2(net227488), .ZN(n404) );
  NAND3_X1 U210 ( .A1(n407), .A2(n406), .A3(n405), .ZN(Y[18]) );
  NAND3_X1 U211 ( .A1(n410), .A2(n409), .A3(n408), .ZN(Y[19]) );
  NAND3_X1 U212 ( .A1(n413), .A2(n412), .A3(n411), .ZN(Y[20]) );
  NAND3_X1 U213 ( .A1(n416), .A2(n415), .A3(n414), .ZN(Y[21]) );
  NAND3_X1 U214 ( .A1(n419), .A2(n418), .A3(n417), .ZN(Y[22]) );
  NAND3_X1 U215 ( .A1(n422), .A2(n421), .A3(n420), .ZN(Y[23]) );
  NAND3_X1 U216 ( .A1(n425), .A2(n424), .A3(n423), .ZN(Y[24]) );
  NAND3_X1 U217 ( .A1(n428), .A2(n427), .A3(n426), .ZN(Y[25]) );
  NAND3_X1 U218 ( .A1(n431), .A2(n430), .A3(n429), .ZN(Y[26]) );
  NAND3_X1 U219 ( .A1(n434), .A2(n433), .A3(n432), .ZN(Y[27]) );
  NAND3_X1 U220 ( .A1(n437), .A2(n436), .A3(n435), .ZN(Y[28]) );
  NAND3_X1 U221 ( .A1(n440), .A2(n439), .A3(n438), .ZN(Y[29]) );
  NAND3_X1 U222 ( .A1(n443), .A2(n442), .A3(n441), .ZN(Y[30]) );
  NAND3_X1 U223 ( .A1(n446), .A2(n445), .A3(n444), .ZN(Y[31]) );
endmodule


module Boothencoder_7 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   net233081, net232889, net227657, net227656, n12, n13, n14, n15, n16,
         n17, n18, n19;
  assign S[2] = net233081;

  CLKBUF_X1 U1 ( .A(n17), .Z(n12) );
  NAND2_X1 U2 ( .A1(n17), .A2(n16), .ZN(n13) );
  INV_X1 U3 ( .A(B[2]), .ZN(n14) );
  AND2_X2 U4 ( .A1(n13), .A2(n14), .ZN(S[0]) );
  BUF_X1 U5 ( .A(B[1]), .Z(n18) );
  AND2_X2 U6 ( .A1(n19), .A2(B[2]), .ZN(net233081) );
  INV_X1 U7 ( .A(n16), .ZN(n15) );
  INV_X1 U8 ( .A(B[1]), .ZN(n16) );
  AND2_X1 U9 ( .A1(n17), .A2(n16), .ZN(n19) );
  INV_X1 U10 ( .A(B[0]), .ZN(n17) );
  BUF_X1 U11 ( .A(n17), .Z(net232889) );
  NAND3_X1 U12 ( .A1(net232889), .A2(n15), .A3(B[2]), .ZN(net227657) );
  XNOR2_X1 U13 ( .A(B[2]), .B(n18), .ZN(net227656) );
  OAI21_X1 U14 ( .B1(net227656), .B2(n12), .A(net227657), .ZN(S[1]) );
endmodule


module mux51_generic_N32_0 ( A, B, C, D, E, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] S;
  output [31:0] Y;
  wire   net227665, net227670, net227687, net227704, net227705, net227762,
         net227798, net227806, net227812, net227814, net227817, net227819,
         net227836, net227841, net232316, net232324, net232322, net233096,
         net233095, net239817, net239882, net240399, net240455, net240475,
         net240474, net241381, net241504, net242000, net242537, net242598,
         net242717, net242036, net232318, net243714, net242004, net239873,
         net227823, net227822, net227821, net227858, net233246, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429;

  BUF_X2 U2 ( .A(net242036), .Z(n303) );
  INV_X1 U3 ( .A(net240475), .ZN(n290) );
  BUF_X1 U4 ( .A(net242036), .Z(net232322) );
  INV_X1 U5 ( .A(net239882), .ZN(n291) );
  BUF_X2 U6 ( .A(S[1]), .Z(net239882) );
  CLKBUF_X1 U7 ( .A(net242598), .Z(n292) );
  NAND2_X1 U8 ( .A1(n296), .A2(n297), .ZN(Y[2]) );
  NAND2_X2 U9 ( .A1(n368), .A2(n304), .ZN(Y[13]) );
  BUF_X1 U10 ( .A(n319), .Z(n293) );
  CLKBUF_X1 U11 ( .A(net242004), .Z(n294) );
  AND2_X2 U12 ( .A1(n308), .A2(net240455), .ZN(net242004) );
  BUF_X2 U13 ( .A(net242004), .Z(net232316) );
  AND2_X2 U14 ( .A1(net227836), .A2(net233096), .ZN(net242717) );
  BUF_X1 U15 ( .A(net242598), .Z(net243714) );
  CLKBUF_X1 U16 ( .A(net240399), .Z(n295) );
  AND2_X1 U17 ( .A1(net227836), .A2(net233096), .ZN(net242598) );
  AND2_X1 U18 ( .A1(n344), .A2(n343), .ZN(n296) );
  NOR2_X1 U19 ( .A1(n341), .A2(n342), .ZN(n297) );
  NAND3_X1 U20 ( .A1(n393), .A2(n392), .A3(n391), .ZN(Y[20]) );
  NAND3_X1 U21 ( .A1(n357), .A2(n359), .A3(n358), .ZN(Y[10]) );
  AND2_X1 U22 ( .A1(n354), .A2(n355), .ZN(n298) );
  AND2_X1 U23 ( .A1(n381), .A2(n379), .ZN(n299) );
  AND3_X1 U24 ( .A1(n331), .A2(n330), .A3(n332), .ZN(n300) );
  AND2_X1 U25 ( .A1(n365), .A2(n364), .ZN(n301) );
  CLKBUF_X3 U26 ( .A(net242036), .Z(n302) );
  BUF_X2 U27 ( .A(S[1]), .Z(n308) );
  AND2_X1 U28 ( .A1(n366), .A2(n367), .ZN(n304) );
  CLKBUF_X1 U29 ( .A(net242036), .Z(net232324) );
  AND2_X1 U30 ( .A1(n310), .A2(S[0]), .ZN(net233096) );
  INV_X1 U31 ( .A(net227670), .ZN(net227687) );
  NOR2_X1 U32 ( .A1(net239882), .A2(net227858), .ZN(n305) );
  AND2_X1 U33 ( .A1(n309), .A2(n310), .ZN(n306) );
  AND2_X1 U34 ( .A1(n309), .A2(n310), .ZN(net240455) );
  AOI22_X1 U35 ( .A1(B[3]), .A2(net242717), .B1(net233246), .B2(E[3]), .ZN(
        n307) );
  NAND4_X1 U36 ( .A1(n307), .A2(net227821), .A3(net227822), .A4(net227823), 
        .ZN(Y[3]) );
  AOI22_X1 U37 ( .A1(E[5]), .A2(net233246), .B1(B[5]), .B2(net242717), .ZN(
        net227812) );
  NAND2_X1 U38 ( .A1(E[4]), .A2(net233246), .ZN(net227817) );
  INV_X1 U39 ( .A(S[1]), .ZN(net227836) );
  NOR2_X1 U40 ( .A1(net239882), .A2(net227858), .ZN(net233246) );
  NOR2_X1 U41 ( .A1(net227858), .A2(n308), .ZN(net242036) );
  AND2_X1 U42 ( .A1(net233095), .A2(n308), .ZN(net239873) );
  NAND2_X1 U43 ( .A1(net241504), .A2(net233095), .ZN(net240474) );
  NAND2_X1 U44 ( .A1(n311), .A2(n309), .ZN(net227858) );
  INV_X1 U45 ( .A(S[0]), .ZN(n309) );
  AND2_X1 U46 ( .A1(n309), .A2(n311), .ZN(net242000) );
  CLKBUF_X1 U47 ( .A(S[2]), .Z(n311) );
  AND2_X1 U48 ( .A1(n310), .A2(S[0]), .ZN(net233095) );
  INV_X1 U49 ( .A(S[2]), .ZN(n310) );
  NAND2_X1 U50 ( .A1(C[3]), .A2(net242004), .ZN(net227823) );
  NAND2_X1 U51 ( .A1(C[5]), .A2(net242004), .ZN(net227814) );
  NAND2_X1 U52 ( .A1(C[7]), .A2(n294), .ZN(net227806) );
  NAND2_X1 U53 ( .A1(C[4]), .A2(net242004), .ZN(net227819) );
  NAND2_X1 U54 ( .A1(A[3]), .A2(net240399), .ZN(net227822) );
  NAND2_X1 U55 ( .A1(net239873), .A2(D[3]), .ZN(net227821) );
  CLKBUF_X1 U56 ( .A(net242004), .Z(net232318) );
  AND2_X2 U57 ( .A1(net227836), .A2(net240455), .ZN(net240399) );
  AND2_X1 U58 ( .A1(net239873), .A2(D[1]), .ZN(net227841) );
  NAND4_X1 U59 ( .A1(n312), .A2(n313), .A3(n314), .A4(n315), .ZN(Y[6]) );
  NAND2_X1 U60 ( .A1(A[6]), .A2(net240399), .ZN(n315) );
  NAND2_X1 U61 ( .A1(C[6]), .A2(n294), .ZN(n314) );
  BUF_X1 U62 ( .A(net232318), .Z(net239817) );
  NAND2_X1 U63 ( .A1(C[15]), .A2(net239817), .ZN(net227762) );
  NAND2_X1 U64 ( .A1(C[9]), .A2(net232318), .ZN(net227798) );
  NAND2_X1 U65 ( .A1(D[6]), .A2(net242537), .ZN(n313) );
  AOI22_X1 U66 ( .A1(E[6]), .A2(net232322), .B1(B[6]), .B2(net243714), .ZN(
        n312) );
  AND2_X1 U67 ( .A1(n308), .A2(net233096), .ZN(net242537) );
  INV_X2 U68 ( .A(net240474), .ZN(net241381) );
  INV_X1 U69 ( .A(net242717), .ZN(net240475) );
  NAND2_X1 U70 ( .A1(n300), .A2(n333), .ZN(Y[0]) );
  NAND2_X1 U71 ( .A1(n338), .A2(n337), .ZN(Y[1]) );
  INV_X1 U72 ( .A(net242537), .ZN(net227670) );
  AND2_X1 U73 ( .A1(n316), .A2(n317), .ZN(n318) );
  NAND2_X1 U74 ( .A1(D[5]), .A2(net242537), .ZN(n316) );
  NAND2_X1 U75 ( .A1(A[5]), .A2(net240399), .ZN(n317) );
  NAND4_X1 U76 ( .A1(n347), .A2(net227817), .A3(n346), .A4(net227819), .ZN(
        Y[4]) );
  CLKBUF_X1 U77 ( .A(n291), .Z(net241504) );
  NAND3_X1 U78 ( .A1(net227762), .A2(n377), .A3(n376), .ZN(Y[15]) );
  NAND2_X2 U79 ( .A1(n380), .A2(n299), .ZN(Y[16]) );
  INV_X1 U80 ( .A(net227665), .ZN(net227704) );
  INV_X1 U81 ( .A(net240399), .ZN(net227665) );
  NAND3_X2 U82 ( .A1(net227798), .A2(n356), .A3(n298), .ZN(Y[9]) );
  NAND3_X1 U83 ( .A1(n360), .A2(n361), .A3(n362), .ZN(Y[11]) );
  NAND3_X1 U84 ( .A1(n318), .A2(net227814), .A3(net227812), .ZN(Y[5]) );
  NAND2_X1 U85 ( .A1(n363), .A2(n301), .ZN(Y[12]) );
  NAND4_X1 U86 ( .A1(n350), .A2(net227806), .A3(n349), .A4(n348), .ZN(Y[7]) );
  NOR2_X1 U87 ( .A1(net227670), .A2(n325), .ZN(n375) );
  INV_X1 U88 ( .A(net227670), .ZN(net227705) );
  NAND2_X1 U89 ( .A1(D[10]), .A2(n423), .ZN(n358) );
  NAND2_X1 U90 ( .A1(E[19]), .A2(n303), .ZN(n389) );
  NAND2_X1 U91 ( .A1(E[21]), .A2(n302), .ZN(n395) );
  NAND2_X1 U92 ( .A1(E[23]), .A2(n302), .ZN(n401) );
  NAND2_X1 U93 ( .A1(E[25]), .A2(n303), .ZN(n408) );
  NAND2_X1 U94 ( .A1(E[27]), .A2(n303), .ZN(n415) );
  NAND2_X1 U95 ( .A1(E[24]), .A2(net232324), .ZN(n405) );
  AOI22_X1 U96 ( .A1(A[24]), .A2(n403), .B1(C[24]), .B2(net232318), .ZN(n404)
         );
  NAND2_X1 U97 ( .A1(E[22]), .A2(n303), .ZN(n398) );
  AOI22_X1 U98 ( .A1(A[22]), .A2(n403), .B1(C[22]), .B2(net232316), .ZN(n397)
         );
  NAND2_X1 U99 ( .A1(E[26]), .A2(n302), .ZN(n411) );
  AOI22_X1 U100 ( .A1(A[26]), .A2(n403), .B1(C[26]), .B2(net239817), .ZN(n410)
         );
  NAND2_X1 U101 ( .A1(E[28]), .A2(n302), .ZN(n418) );
  AOI22_X1 U102 ( .A1(A[28]), .A2(n403), .B1(C[28]), .B2(net232318), .ZN(n417)
         );
  NAND2_X1 U103 ( .A1(E[20]), .A2(n302), .ZN(n392) );
  NAND3_X1 U104 ( .A1(n387), .A2(n386), .A3(n385), .ZN(Y[18]) );
  NAND2_X1 U105 ( .A1(E[18]), .A2(n303), .ZN(n386) );
  NAND3_X1 U106 ( .A1(n373), .A2(n372), .A3(n371), .ZN(Y[14]) );
  NAND2_X1 U107 ( .A1(D[11]), .A2(n413), .ZN(n361) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(net227687), .ZN(n364) );
  NAND2_X1 U109 ( .A1(E[17]), .A2(net232324), .ZN(n383) );
  AOI21_X1 U110 ( .B1(E[16]), .B2(n302), .A(n378), .ZN(n381) );
  NAND2_X1 U111 ( .A1(E[29]), .A2(n303), .ZN(n421) );
  NAND2_X1 U112 ( .A1(E[30]), .A2(n302), .ZN(n425) );
  NAND2_X1 U113 ( .A1(E[31]), .A2(net232324), .ZN(n428) );
  AOI22_X1 U114 ( .A1(A[31]), .A2(n295), .B1(C[31]), .B2(net232316), .ZN(n427)
         );
  NAND2_X1 U115 ( .A1(D[13]), .A2(net227705), .ZN(n367) );
  AOI22_X1 U116 ( .A1(A[27]), .A2(net227704), .B1(C[27]), .B2(net232316), .ZN(
        n414) );
  AOI22_X1 U117 ( .A1(A[25]), .A2(net227704), .B1(C[25]), .B2(net232316), .ZN(
        n407) );
  AOI22_X1 U118 ( .A1(A[23]), .A2(net227704), .B1(C[23]), .B2(net232316), .ZN(
        n400) );
  NAND2_X1 U119 ( .A1(net227836), .A2(n306), .ZN(n319) );
  INV_X1 U120 ( .A(n320), .ZN(n423) );
  INV_X1 U121 ( .A(n320), .ZN(n413) );
  NOR2_X1 U122 ( .A1(n320), .A2(n324), .ZN(n370) );
  NAND3_X2 U123 ( .A1(n351), .A2(n352), .A3(n353), .ZN(Y[8]) );
  AOI22_X1 U124 ( .A1(A[11]), .A2(n403), .B1(C[11]), .B2(net232318), .ZN(n362)
         );
  NAND2_X1 U125 ( .A1(C[16]), .A2(net239817), .ZN(n380) );
  INV_X1 U126 ( .A(n293), .ZN(n403) );
  NOR2_X1 U127 ( .A1(n339), .A2(n319), .ZN(n342) );
  AOI22_X1 U128 ( .A1(A[21]), .A2(net227704), .B1(C[21]), .B2(net232318), .ZN(
        n394) );
  AOI22_X1 U129 ( .A1(A[17]), .A2(net227704), .B1(C[17]), .B2(net239817), .ZN(
        n382) );
  AOI22_X1 U130 ( .A1(A[20]), .A2(n403), .B1(C[20]), .B2(net232318), .ZN(n391)
         );
  AOI22_X1 U131 ( .A1(A[19]), .A2(net227704), .B1(C[19]), .B2(net232316), .ZN(
        n388) );
  AOI22_X1 U132 ( .A1(A[18]), .A2(n403), .B1(C[18]), .B2(net232316), .ZN(n385)
         );
  AOI22_X1 U133 ( .A1(C[10]), .A2(net232316), .B1(A[10]), .B2(net240399), .ZN(
        n357) );
  NOR2_X1 U134 ( .A1(net240474), .A2(n322), .ZN(n378) );
  NOR2_X1 U135 ( .A1(net240475), .A2(n326), .ZN(n369) );
  NOR2_X1 U136 ( .A1(net240474), .A2(n321), .ZN(n374) );
  AOI211_X1 U137 ( .C1(E[14]), .C2(n302), .A(n370), .B(n369), .ZN(n371) );
  NAND2_X1 U138 ( .A1(E[8]), .A2(n302), .ZN(n352) );
  NAND2_X1 U139 ( .A1(net239882), .A2(net233095), .ZN(n320) );
  AOI22_X1 U140 ( .A1(A[30]), .A2(n403), .B1(C[30]), .B2(net232316), .ZN(n424)
         );
  AOI22_X1 U141 ( .A1(A[29]), .A2(net227704), .B1(C[29]), .B2(net232316), .ZN(
        n420) );
  NAND2_X1 U142 ( .A1(C[14]), .A2(net239817), .ZN(n373) );
  AOI22_X1 U143 ( .A1(D[31]), .A2(net227687), .B1(B[31]), .B2(net241381), .ZN(
        n429) );
  AOI22_X1 U144 ( .A1(D[28]), .A2(net227687), .B1(B[28]), .B2(net241381), .ZN(
        n419) );
  AOI22_X1 U145 ( .A1(D[21]), .A2(n413), .B1(B[21]), .B2(net241381), .ZN(n396)
         );
  AOI22_X1 U146 ( .A1(D[20]), .A2(net227687), .B1(B[20]), .B2(net241381), .ZN(
        n393) );
  AOI22_X1 U147 ( .A1(D[17]), .A2(n423), .B1(B[17]), .B2(net241381), .ZN(n384)
         );
  AOI22_X1 U148 ( .A1(D[19]), .A2(net227687), .B1(B[19]), .B2(net241381), .ZN(
        n390) );
  AOI22_X1 U149 ( .A1(D[18]), .A2(n423), .B1(B[18]), .B2(net241381), .ZN(n387)
         );
  AOI22_X1 U150 ( .A1(A[12]), .A2(net240399), .B1(B[12]), .B2(net242717), .ZN(
        n365) );
  AOI22_X1 U151 ( .A1(C[8]), .A2(net232316), .B1(B[8]), .B2(net242717), .ZN(
        n353) );
  AOI22_X1 U152 ( .A1(E[9]), .A2(n302), .B1(B[9]), .B2(net242717), .ZN(n356)
         );
  AOI22_X1 U153 ( .A1(C[12]), .A2(net232316), .B1(E[12]), .B2(net232324), .ZN(
        n363) );
  AOI211_X1 U154 ( .C1(E[15]), .C2(n303), .A(n375), .B(n374), .ZN(n376) );
  NAND2_X1 U155 ( .A1(n306), .A2(n308), .ZN(n345) );
  AOI22_X1 U156 ( .A1(D[30]), .A2(n423), .B1(B[30]), .B2(net241381), .ZN(n426)
         );
  AOI22_X1 U157 ( .A1(D[29]), .A2(net227687), .B1(B[29]), .B2(net241381), .ZN(
        n422) );
  AOI22_X1 U158 ( .A1(D[27]), .A2(n413), .B1(B[27]), .B2(net241381), .ZN(n416)
         );
  AOI22_X1 U159 ( .A1(D[26]), .A2(net227687), .B1(B[26]), .B2(net241381), .ZN(
        n412) );
  AOI22_X1 U160 ( .A1(D[25]), .A2(net227705), .B1(B[25]), .B2(net241381), .ZN(
        n409) );
  AOI22_X1 U161 ( .A1(D[24]), .A2(n413), .B1(B[24]), .B2(net241381), .ZN(n406)
         );
  AOI22_X1 U162 ( .A1(D[23]), .A2(net227687), .B1(B[23]), .B2(n292), .ZN(n402)
         );
  AOI22_X1 U163 ( .A1(D[22]), .A2(net227687), .B1(B[22]), .B2(n290), .ZN(n399)
         );
  AOI22_X1 U164 ( .A1(B[13]), .A2(n292), .B1(E[13]), .B2(n302), .ZN(n366) );
  AOI22_X1 U165 ( .A1(B[10]), .A2(n292), .B1(E[10]), .B2(n303), .ZN(n359) );
  AOI22_X1 U166 ( .A1(B[11]), .A2(n292), .B1(E[11]), .B2(n303), .ZN(n360) );
  AOI22_X1 U167 ( .A1(A[13]), .A2(n403), .B1(C[13]), .B2(net239817), .ZN(n368)
         );
  INV_X1 U168 ( .A(B[15]), .ZN(n321) );
  INV_X1 U169 ( .A(B[16]), .ZN(n322) );
  INV_X1 U170 ( .A(B[0]), .ZN(n323) );
  INV_X1 U171 ( .A(D[14]), .ZN(n324) );
  INV_X1 U172 ( .A(D[15]), .ZN(n325) );
  INV_X1 U173 ( .A(B[14]), .ZN(n326) );
  INV_X1 U174 ( .A(E[0]), .ZN(n327) );
  NOR2_X1 U175 ( .A1(n327), .A2(net239882), .ZN(n329) );
  NOR2_X1 U176 ( .A1(n323), .A2(net239882), .ZN(n328) );
  AOI22_X1 U177 ( .A1(net242000), .A2(n329), .B1(n328), .B2(net233095), .ZN(
        n333) );
  NAND3_X1 U178 ( .A1(net239882), .A2(D[0]), .A3(net233095), .ZN(n332) );
  NAND3_X1 U179 ( .A1(net239882), .A2(C[0]), .A3(n306), .ZN(n331) );
  NAND3_X1 U180 ( .A1(net227836), .A2(A[0]), .A3(n306), .ZN(n330) );
  INV_X1 U181 ( .A(C[1]), .ZN(n335) );
  INV_X1 U182 ( .A(A[1]), .ZN(n334) );
  OAI22_X1 U183 ( .A1(n345), .A2(n335), .B1(n319), .B2(n334), .ZN(n336) );
  NOR2_X1 U184 ( .A1(n336), .A2(net227841), .ZN(n338) );
  AOI22_X1 U185 ( .A1(n305), .A2(E[1]), .B1(B[1]), .B2(net242717), .ZN(n337)
         );
  AOI22_X1 U186 ( .A1(n305), .A2(E[2]), .B1(net242598), .B2(B[2]), .ZN(n344)
         );
  NAND2_X1 U187 ( .A1(D[2]), .A2(net242537), .ZN(n343) );
  INV_X1 U188 ( .A(A[2]), .ZN(n339) );
  INV_X1 U189 ( .A(C[2]), .ZN(n340) );
  NOR2_X1 U190 ( .A1(n345), .A2(n340), .ZN(n341) );
  NAND2_X1 U191 ( .A1(D[4]), .A2(net242537), .ZN(n347) );
  AOI22_X1 U192 ( .A1(A[4]), .A2(net240399), .B1(B[4]), .B2(net242598), .ZN(
        n346) );
  AOI22_X1 U193 ( .A1(E[7]), .A2(net232322), .B1(B[7]), .B2(net243714), .ZN(
        n350) );
  NAND2_X1 U194 ( .A1(D[7]), .A2(n413), .ZN(n349) );
  NAND2_X1 U195 ( .A1(A[7]), .A2(net240399), .ZN(n348) );
  AOI22_X1 U196 ( .A1(A[8]), .A2(net240399), .B1(D[8]), .B2(net227705), .ZN(
        n351) );
  NAND2_X1 U197 ( .A1(D[9]), .A2(n423), .ZN(n355) );
  NAND2_X1 U198 ( .A1(A[9]), .A2(net240399), .ZN(n354) );
  NAND2_X1 U199 ( .A1(A[14]), .A2(n295), .ZN(n372) );
  NAND2_X1 U200 ( .A1(A[15]), .A2(n295), .ZN(n377) );
  AOI22_X1 U201 ( .A1(A[16]), .A2(net227704), .B1(D[16]), .B2(net227687), .ZN(
        n379) );
  NAND3_X1 U202 ( .A1(n384), .A2(n383), .A3(n382), .ZN(Y[17]) );
  NAND3_X1 U203 ( .A1(n390), .A2(n389), .A3(n388), .ZN(Y[19]) );
  NAND3_X1 U204 ( .A1(n396), .A2(n395), .A3(n394), .ZN(Y[21]) );
  NAND3_X1 U205 ( .A1(n399), .A2(n398), .A3(n397), .ZN(Y[22]) );
  NAND3_X1 U206 ( .A1(n402), .A2(n401), .A3(n400), .ZN(Y[23]) );
  NAND3_X1 U207 ( .A1(n406), .A2(n405), .A3(n404), .ZN(Y[24]) );
  NAND3_X1 U208 ( .A1(n409), .A2(n408), .A3(n407), .ZN(Y[25]) );
  NAND3_X1 U209 ( .A1(n412), .A2(n411), .A3(n410), .ZN(Y[26]) );
  NAND3_X1 U210 ( .A1(n416), .A2(n415), .A3(n414), .ZN(Y[27]) );
  NAND3_X1 U211 ( .A1(n419), .A2(n418), .A3(n417), .ZN(Y[28]) );
  NAND3_X1 U212 ( .A1(n422), .A2(n421), .A3(n420), .ZN(Y[29]) );
  NAND3_X1 U213 ( .A1(n426), .A2(n425), .A3(n424), .ZN(Y[30]) );
  NAND3_X1 U214 ( .A1(n429), .A2(n428), .A3(n427), .ZN(Y[31]) );
endmodule


module Boothencoder_0 ( B, S );
  input [2:0] B;
  output [2:0] S;
  wire   net227859, net242606, n11, n12, n13, n14, n15, n16;

  NAND2_X1 U1 ( .A1(n15), .A2(n11), .ZN(n12) );
  AND2_X1 U2 ( .A1(B[0]), .A2(B[1]), .ZN(n11) );
  OAI21_X1 U3 ( .B1(n14), .B2(n15), .A(n12), .ZN(S[1]) );
  INV_X1 U4 ( .A(B[1]), .ZN(n16) );
  INV_X1 U5 ( .A(n16), .ZN(net242606) );
  AOI21_X1 U6 ( .B1(n16), .B2(n13), .A(B[2]), .ZN(S[0]) );
  INV_X1 U7 ( .A(B[2]), .ZN(n15) );
  INV_X1 U8 ( .A(B[0]), .ZN(n13) );
  XNOR2_X1 U9 ( .A(B[1]), .B(B[0]), .ZN(n14) );
  NAND2_X1 U10 ( .A1(B[2]), .A2(n13), .ZN(net227859) );
  NOR2_X1 U11 ( .A1(net227859), .A2(net242606), .ZN(S[2]) );
endmodule


module SHIFTER_GENERIC_N32_DW_rbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \MR_int[1][31] , \MR_int[1][30] , \MR_int[1][29] , \MR_int[1][28] ,
         \MR_int[1][27] , \MR_int[1][26] , \MR_int[1][25] , \MR_int[1][24] ,
         \MR_int[1][23] , \MR_int[1][22] , \MR_int[1][21] , \MR_int[1][20] ,
         \MR_int[1][19] , \MR_int[1][18] , \MR_int[1][17] , \MR_int[1][16] ,
         \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] , \MR_int[1][12] ,
         \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] , \MR_int[1][8] ,
         \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] , \MR_int[1][4] ,
         \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] , \MR_int[1][0] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][28] ,
         \MR_int[2][27] , \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] ,
         \MR_int[2][23] , \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] ,
         \MR_int[2][19] , \MR_int[2][18] , \MR_int[2][17] , \MR_int[2][16] ,
         \MR_int[2][15] , \MR_int[2][14] , \MR_int[2][13] , \MR_int[2][12] ,
         \MR_int[2][11] , \MR_int[2][10] , \MR_int[2][9] , \MR_int[2][8] ,
         \MR_int[2][7] , \MR_int[2][6] , \MR_int[2][5] , \MR_int[2][4] ,
         \MR_int[2][3] , \MR_int[2][2] , \MR_int[2][1] , \MR_int[2][0] ,
         \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] , \MR_int[3][28] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][22] , \MR_int[3][21] , \MR_int[3][20] ,
         \MR_int[3][19] , \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] ,
         \MR_int[3][15] , \MR_int[3][14] , \MR_int[3][13] , \MR_int[3][12] ,
         \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] , \MR_int[3][8] ,
         \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][5] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[3][0] ,
         \MR_int[4][31] , \MR_int[4][30] , \MR_int[4][29] , \MR_int[4][28] ,
         \MR_int[4][27] , \MR_int[4][26] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][23] , \MR_int[4][22] , \MR_int[4][21] , \MR_int[4][20] ,
         \MR_int[4][19] , \MR_int[4][18] , \MR_int[4][17] , \MR_int[4][16] ,
         \MR_int[4][15] , \MR_int[4][14] , \MR_int[4][13] , \MR_int[4][12] ,
         \MR_int[4][11] , \MR_int[4][10] , \MR_int[4][9] , \MR_int[4][8] ,
         \MR_int[4][7] , \MR_int[4][6] , \MR_int[4][5] , \MR_int[4][4] ,
         \MR_int[4][3] , \MR_int[4][2] , \MR_int[4][1] , \MR_int[4][0] , n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;

  MUX2_X1 M1_4_31 ( .A(\MR_int[4][31] ), .B(\MR_int[4][15] ), .S(n18), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\MR_int[4][30] ), .B(\MR_int[4][14] ), .S(n18), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\MR_int[4][29] ), .B(\MR_int[4][13] ), .S(n18), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\MR_int[4][28] ), .B(\MR_int[4][12] ), .S(n18), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\MR_int[4][27] ), .B(\MR_int[4][11] ), .S(n18), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\MR_int[4][26] ), .B(\MR_int[4][10] ), .S(n18), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\MR_int[4][25] ), .B(\MR_int[4][9] ), .S(n18), .Z(B[25]) );
  MUX2_X1 M1_4_24 ( .A(\MR_int[4][24] ), .B(\MR_int[4][8] ), .S(n18), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\MR_int[4][23] ), .B(\MR_int[4][7] ), .S(n17), .Z(B[23]) );
  MUX2_X1 M1_4_22 ( .A(\MR_int[4][22] ), .B(\MR_int[4][6] ), .S(n17), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\MR_int[4][21] ), .B(\MR_int[4][5] ), .S(n17), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\MR_int[4][20] ), .B(\MR_int[4][4] ), .S(n17), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\MR_int[4][19] ), .B(\MR_int[4][3] ), .S(n17), .Z(B[19]) );
  MUX2_X1 M1_4_18 ( .A(\MR_int[4][18] ), .B(\MR_int[4][2] ), .S(n17), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\MR_int[4][17] ), .B(\MR_int[4][1] ), .S(n17), .Z(B[17]) );
  MUX2_X1 M1_4_16 ( .A(\MR_int[4][16] ), .B(\MR_int[4][0] ), .S(n17), .Z(B[16]) );
  MUX2_X1 M1_4_15 ( .A(\MR_int[4][15] ), .B(\MR_int[4][31] ), .S(n17), .Z(
        B[15]) );
  MUX2_X1 M1_4_14 ( .A(\MR_int[4][14] ), .B(\MR_int[4][30] ), .S(n17), .Z(
        B[14]) );
  MUX2_X1 M1_4_13 ( .A(\MR_int[4][13] ), .B(\MR_int[4][29] ), .S(n17), .Z(
        B[13]) );
  MUX2_X1 M1_4_12 ( .A(\MR_int[4][12] ), .B(\MR_int[4][28] ), .S(n17), .Z(
        B[12]) );
  MUX2_X1 M1_4_11 ( .A(\MR_int[4][11] ), .B(\MR_int[4][27] ), .S(n16), .Z(
        B[11]) );
  MUX2_X1 M1_4_10 ( .A(\MR_int[4][10] ), .B(\MR_int[4][26] ), .S(n16), .Z(
        B[10]) );
  MUX2_X1 M1_4_9 ( .A(\MR_int[4][9] ), .B(\MR_int[4][25] ), .S(n16), .Z(B[9])
         );
  MUX2_X1 M1_4_8 ( .A(\MR_int[4][8] ), .B(\MR_int[4][24] ), .S(n16), .Z(B[8])
         );
  MUX2_X1 M1_4_7 ( .A(\MR_int[4][7] ), .B(\MR_int[4][23] ), .S(n16), .Z(B[7])
         );
  MUX2_X1 M1_4_6 ( .A(\MR_int[4][6] ), .B(\MR_int[4][22] ), .S(n16), .Z(B[6])
         );
  MUX2_X1 M1_4_5 ( .A(\MR_int[4][5] ), .B(\MR_int[4][21] ), .S(n16), .Z(B[5])
         );
  MUX2_X1 M1_4_4 ( .A(\MR_int[4][4] ), .B(\MR_int[4][20] ), .S(n16), .Z(B[4])
         );
  MUX2_X1 M1_4_3 ( .A(\MR_int[4][3] ), .B(\MR_int[4][19] ), .S(n16), .Z(B[3])
         );
  MUX2_X1 M1_4_2 ( .A(\MR_int[4][2] ), .B(\MR_int[4][18] ), .S(n16), .Z(B[2])
         );
  MUX2_X1 M1_4_1 ( .A(\MR_int[4][1] ), .B(\MR_int[4][17] ), .S(n16), .Z(B[1])
         );
  MUX2_X1 M1_4_0 ( .A(\MR_int[4][0] ), .B(\MR_int[4][16] ), .S(n16), .Z(B[0])
         );
  MUX2_X1 M1_3_31_0 ( .A(\MR_int[3][31] ), .B(\MR_int[3][7] ), .S(n27), .Z(
        \MR_int[4][31] ) );
  MUX2_X1 M1_3_30_0 ( .A(\MR_int[3][30] ), .B(\MR_int[3][6] ), .S(n27), .Z(
        \MR_int[4][30] ) );
  MUX2_X1 M1_3_29_0 ( .A(\MR_int[3][29] ), .B(\MR_int[3][5] ), .S(n27), .Z(
        \MR_int[4][29] ) );
  MUX2_X1 M1_3_28_0 ( .A(\MR_int[3][28] ), .B(\MR_int[3][4] ), .S(n27), .Z(
        \MR_int[4][28] ) );
  MUX2_X1 M1_3_27_0 ( .A(\MR_int[3][27] ), .B(\MR_int[3][3] ), .S(n27), .Z(
        \MR_int[4][27] ) );
  MUX2_X1 M1_3_26_0 ( .A(\MR_int[3][26] ), .B(\MR_int[3][2] ), .S(n27), .Z(
        \MR_int[4][26] ) );
  MUX2_X1 M1_3_25_0 ( .A(\MR_int[3][25] ), .B(\MR_int[3][1] ), .S(n27), .Z(
        \MR_int[4][25] ) );
  MUX2_X1 M1_3_24_0 ( .A(\MR_int[3][24] ), .B(\MR_int[3][0] ), .S(n27), .Z(
        \MR_int[4][24] ) );
  MUX2_X1 M1_3_23_0 ( .A(\MR_int[3][23] ), .B(\MR_int[3][31] ), .S(n26), .Z(
        \MR_int[4][23] ) );
  MUX2_X1 M1_3_22_0 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(n26), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_21_0 ( .A(\MR_int[3][21] ), .B(\MR_int[3][29] ), .S(n26), .Z(
        \MR_int[4][21] ) );
  MUX2_X1 M1_3_20_0 ( .A(\MR_int[3][20] ), .B(\MR_int[3][28] ), .S(n26), .Z(
        \MR_int[4][20] ) );
  MUX2_X1 M1_3_19_0 ( .A(\MR_int[3][19] ), .B(\MR_int[3][27] ), .S(n26), .Z(
        \MR_int[4][19] ) );
  MUX2_X1 M1_3_18_0 ( .A(\MR_int[3][18] ), .B(\MR_int[3][26] ), .S(n26), .Z(
        \MR_int[4][18] ) );
  MUX2_X1 M1_3_17_0 ( .A(\MR_int[3][17] ), .B(\MR_int[3][25] ), .S(n26), .Z(
        \MR_int[4][17] ) );
  MUX2_X1 M1_3_16_0 ( .A(\MR_int[3][16] ), .B(\MR_int[3][24] ), .S(n26), .Z(
        \MR_int[4][16] ) );
  MUX2_X1 M1_3_15_0 ( .A(\MR_int[3][15] ), .B(\MR_int[3][23] ), .S(n26), .Z(
        \MR_int[4][15] ) );
  MUX2_X1 M1_3_14_0 ( .A(\MR_int[3][14] ), .B(\MR_int[3][22] ), .S(n26), .Z(
        \MR_int[4][14] ) );
  MUX2_X1 M1_3_13_0 ( .A(\MR_int[3][13] ), .B(\MR_int[3][21] ), .S(n26), .Z(
        \MR_int[4][13] ) );
  MUX2_X1 M1_3_12_0 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(n26), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(n25), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_10_0 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(n25), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 M1_3_9_0 ( .A(\MR_int[3][9] ), .B(\MR_int[3][17] ), .S(n25), .Z(
        \MR_int[4][9] ) );
  MUX2_X1 M1_3_8_0 ( .A(\MR_int[3][8] ), .B(\MR_int[3][16] ), .S(n25), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 M1_3_7 ( .A(\MR_int[3][7] ), .B(\MR_int[3][15] ), .S(n25), .Z(
        \MR_int[4][7] ) );
  MUX2_X1 M1_3_6 ( .A(\MR_int[3][6] ), .B(\MR_int[3][14] ), .S(n25), .Z(
        \MR_int[4][6] ) );
  MUX2_X1 M1_3_5 ( .A(\MR_int[3][5] ), .B(\MR_int[3][13] ), .S(n25), .Z(
        \MR_int[4][5] ) );
  MUX2_X1 M1_3_4 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(n25), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(n25), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(n25), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_3_1 ( .A(\MR_int[3][1] ), .B(\MR_int[3][9] ), .S(n25), .Z(
        \MR_int[4][1] ) );
  MUX2_X1 M1_3_0 ( .A(\MR_int[3][0] ), .B(\MR_int[3][8] ), .S(n25), .Z(
        \MR_int[4][0] ) );
  MUX2_X1 M1_2_31_0 ( .A(\MR_int[2][31] ), .B(\MR_int[2][3] ), .S(n24), .Z(
        \MR_int[3][31] ) );
  MUX2_X1 M1_2_30_0 ( .A(\MR_int[2][30] ), .B(\MR_int[2][2] ), .S(n24), .Z(
        \MR_int[3][30] ) );
  MUX2_X1 M1_2_29_0 ( .A(\MR_int[2][29] ), .B(\MR_int[2][1] ), .S(n24), .Z(
        \MR_int[3][29] ) );
  MUX2_X1 M1_2_28_0 ( .A(\MR_int[2][28] ), .B(\MR_int[2][0] ), .S(n24), .Z(
        \MR_int[3][28] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n24), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 M1_2_26_0 ( .A(\MR_int[2][26] ), .B(\MR_int[2][30] ), .S(n24), .Z(
        \MR_int[3][26] ) );
  MUX2_X1 M1_2_25_0 ( .A(\MR_int[2][25] ), .B(\MR_int[2][29] ), .S(n24), .Z(
        \MR_int[3][25] ) );
  MUX2_X1 M1_2_24_0 ( .A(\MR_int[2][24] ), .B(\MR_int[2][28] ), .S(n24), .Z(
        \MR_int[3][24] ) );
  MUX2_X1 M1_2_23_0 ( .A(\MR_int[2][23] ), .B(\MR_int[2][27] ), .S(n23), .Z(
        \MR_int[3][23] ) );
  MUX2_X1 M1_2_22_0 ( .A(\MR_int[2][22] ), .B(\MR_int[2][26] ), .S(n23), .Z(
        \MR_int[3][22] ) );
  MUX2_X1 M1_2_21_0 ( .A(\MR_int[2][21] ), .B(\MR_int[2][25] ), .S(n23), .Z(
        \MR_int[3][21] ) );
  MUX2_X1 M1_2_20_0 ( .A(\MR_int[2][20] ), .B(\MR_int[2][24] ), .S(n23), .Z(
        \MR_int[3][20] ) );
  MUX2_X1 M1_2_19_0 ( .A(\MR_int[2][19] ), .B(\MR_int[2][23] ), .S(n23), .Z(
        \MR_int[3][19] ) );
  MUX2_X1 M1_2_18_0 ( .A(\MR_int[2][18] ), .B(\MR_int[2][22] ), .S(n23), .Z(
        \MR_int[3][18] ) );
  MUX2_X1 M1_2_17_0 ( .A(\MR_int[2][17] ), .B(\MR_int[2][21] ), .S(n23), .Z(
        \MR_int[3][17] ) );
  MUX2_X1 M1_2_16_0 ( .A(\MR_int[2][16] ), .B(\MR_int[2][20] ), .S(n23), .Z(
        \MR_int[3][16] ) );
  MUX2_X1 M1_2_15_0 ( .A(\MR_int[2][15] ), .B(\MR_int[2][19] ), .S(n23), .Z(
        \MR_int[3][15] ) );
  MUX2_X1 M1_2_14_0 ( .A(\MR_int[2][14] ), .B(\MR_int[2][18] ), .S(n23), .Z(
        \MR_int[3][14] ) );
  MUX2_X1 M1_2_13_0 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(n23), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 M1_2_12_0 ( .A(\MR_int[2][12] ), .B(\MR_int[2][16] ), .S(n23), .Z(
        \MR_int[3][12] ) );
  MUX2_X1 M1_2_11_0 ( .A(\MR_int[2][11] ), .B(\MR_int[2][15] ), .S(n22), .Z(
        \MR_int[3][11] ) );
  MUX2_X1 M1_2_10_0 ( .A(\MR_int[2][10] ), .B(\MR_int[2][14] ), .S(n22), .Z(
        \MR_int[3][10] ) );
  MUX2_X1 M1_2_9_0 ( .A(\MR_int[2][9] ), .B(\MR_int[2][13] ), .S(n22), .Z(
        \MR_int[3][9] ) );
  MUX2_X1 M1_2_8_0 ( .A(\MR_int[2][8] ), .B(\MR_int[2][12] ), .S(n22), .Z(
        \MR_int[3][8] ) );
  MUX2_X1 M1_2_7_0 ( .A(\MR_int[2][7] ), .B(\MR_int[2][11] ), .S(n22), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(n22), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(n22), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(n22), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(n22), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_2_2 ( .A(\MR_int[2][2] ), .B(\MR_int[2][6] ), .S(n22), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 M1_2_1 ( .A(\MR_int[2][1] ), .B(\MR_int[2][5] ), .S(n22), .Z(
        \MR_int[3][1] ) );
  MUX2_X1 M1_2_0 ( .A(\MR_int[2][0] ), .B(\MR_int[2][4] ), .S(n22), .Z(
        \MR_int[3][0] ) );
  MUX2_X1 M1_1_31_0 ( .A(\MR_int[1][31] ), .B(\MR_int[1][1] ), .S(n21), .Z(
        \MR_int[2][31] ) );
  MUX2_X1 M1_1_30_0 ( .A(\MR_int[1][30] ), .B(\MR_int[1][0] ), .S(n21), .Z(
        \MR_int[2][30] ) );
  MUX2_X1 M1_1_29_0 ( .A(\MR_int[1][29] ), .B(\MR_int[1][31] ), .S(n21), .Z(
        \MR_int[2][29] ) );
  MUX2_X1 M1_1_28_0 ( .A(\MR_int[1][28] ), .B(\MR_int[1][30] ), .S(n21), .Z(
        \MR_int[2][28] ) );
  MUX2_X1 M1_1_27_0 ( .A(\MR_int[1][27] ), .B(\MR_int[1][29] ), .S(n21), .Z(
        \MR_int[2][27] ) );
  MUX2_X1 M1_1_26_0 ( .A(\MR_int[1][26] ), .B(\MR_int[1][28] ), .S(n21), .Z(
        \MR_int[2][26] ) );
  MUX2_X1 M1_1_25_0 ( .A(\MR_int[1][25] ), .B(\MR_int[1][27] ), .S(n21), .Z(
        \MR_int[2][25] ) );
  MUX2_X1 M1_1_24_0 ( .A(\MR_int[1][24] ), .B(\MR_int[1][26] ), .S(n21), .Z(
        \MR_int[2][24] ) );
  MUX2_X1 M1_1_23_0 ( .A(\MR_int[1][23] ), .B(\MR_int[1][25] ), .S(n20), .Z(
        \MR_int[2][23] ) );
  MUX2_X1 M1_1_22_0 ( .A(\MR_int[1][22] ), .B(\MR_int[1][24] ), .S(n20), .Z(
        \MR_int[2][22] ) );
  MUX2_X1 M1_1_21_0 ( .A(\MR_int[1][21] ), .B(\MR_int[1][23] ), .S(n20), .Z(
        \MR_int[2][21] ) );
  MUX2_X1 M1_1_20_0 ( .A(\MR_int[1][20] ), .B(\MR_int[1][22] ), .S(n20), .Z(
        \MR_int[2][20] ) );
  MUX2_X1 M1_1_19_0 ( .A(\MR_int[1][19] ), .B(\MR_int[1][21] ), .S(n20), .Z(
        \MR_int[2][19] ) );
  MUX2_X1 M1_1_18_0 ( .A(\MR_int[1][18] ), .B(\MR_int[1][20] ), .S(n20), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 M1_1_17_0 ( .A(\MR_int[1][17] ), .B(\MR_int[1][19] ), .S(n20), .Z(
        \MR_int[2][17] ) );
  MUX2_X1 M1_1_16_0 ( .A(\MR_int[1][16] ), .B(\MR_int[1][18] ), .S(n20), .Z(
        \MR_int[2][16] ) );
  MUX2_X1 M1_1_15_0 ( .A(\MR_int[1][15] ), .B(\MR_int[1][17] ), .S(n20), .Z(
        \MR_int[2][15] ) );
  MUX2_X1 M1_1_14_0 ( .A(\MR_int[1][14] ), .B(\MR_int[1][16] ), .S(n20), .Z(
        \MR_int[2][14] ) );
  MUX2_X1 M1_1_13_0 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(n20), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 M1_1_12_0 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(n20), .Z(
        \MR_int[2][12] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(n19), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(n19), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_9_0 ( .A(\MR_int[1][9] ), .B(\MR_int[1][11] ), .S(n19), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 M1_1_8_0 ( .A(\MR_int[1][8] ), .B(\MR_int[1][10] ), .S(n19), .Z(
        \MR_int[2][8] ) );
  MUX2_X1 M1_1_7_0 ( .A(\MR_int[1][7] ), .B(\MR_int[1][9] ), .S(n19), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 M1_1_6_0 ( .A(\MR_int[1][6] ), .B(\MR_int[1][8] ), .S(n19), .Z(
        \MR_int[2][6] ) );
  MUX2_X1 M1_1_5_0 ( .A(\MR_int[1][5] ), .B(\MR_int[1][7] ), .S(n19), .Z(
        \MR_int[2][5] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(n19), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(n19), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_2_0 ( .A(\MR_int[1][2] ), .B(\MR_int[1][4] ), .S(n19), .Z(
        \MR_int[2][2] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\MR_int[1][3] ), .S(n19), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_1_0 ( .A(\MR_int[1][0] ), .B(\MR_int[1][2] ), .S(n19), .Z(
        \MR_int[2][0] ) );
  MUX2_X1 M1_0_31_0 ( .A(A[31]), .B(A[0]), .S(SH[0]), .Z(\MR_int[1][31] ) );
  MUX2_X1 M1_0_30_0 ( .A(A[30]), .B(A[31]), .S(SH[0]), .Z(\MR_int[1][30] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(SH[0]), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(SH[0]), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_27_0 ( .A(A[27]), .B(A[28]), .S(SH[0]), .Z(\MR_int[1][27] ) );
  MUX2_X1 M1_0_26_0 ( .A(A[26]), .B(A[27]), .S(SH[0]), .Z(\MR_int[1][26] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(SH[0]), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(SH[0]), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_23_0 ( .A(A[23]), .B(A[24]), .S(SH[0]), .Z(\MR_int[1][23] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(SH[0]), .Z(\MR_int[1][22] ) );
  MUX2_X1 M1_0_21_0 ( .A(A[21]), .B(A[22]), .S(SH[0]), .Z(\MR_int[1][21] ) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(SH[0]), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_19_0 ( .A(A[19]), .B(A[20]), .S(SH[0]), .Z(\MR_int[1][19] ) );
  MUX2_X1 M1_0_18_0 ( .A(A[18]), .B(A[19]), .S(SH[0]), .Z(\MR_int[1][18] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(SH[0]), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(SH[0]), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_15_0 ( .A(A[15]), .B(A[16]), .S(SH[0]), .Z(\MR_int[1][15] ) );
  MUX2_X1 M1_0_14_0 ( .A(A[14]), .B(A[15]), .S(SH[0]), .Z(\MR_int[1][14] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(SH[0]), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_12_0 ( .A(A[12]), .B(A[13]), .S(SH[0]), .Z(\MR_int[1][12] ) );
  MUX2_X1 M1_0_11_0 ( .A(A[11]), .B(A[12]), .S(SH[0]), .Z(\MR_int[1][11] ) );
  MUX2_X1 M1_0_10_0 ( .A(A[10]), .B(A[11]), .S(SH[0]), .Z(\MR_int[1][10] ) );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(SH[0]), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(SH[0]), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_7_0 ( .A(A[7]), .B(A[8]), .S(SH[0]), .Z(\MR_int[1][7] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(SH[0]), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(SH[0]), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(SH[0]), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_3_0 ( .A(A[3]), .B(A[4]), .S(SH[0]), .Z(\MR_int[1][3] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(SH[0]), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(SH[0]), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_0_0 ( .A(A[0]), .B(A[1]), .S(SH[0]), .Z(\MR_int[1][0] ) );
  CLKBUF_X1 U2 ( .A(SH[3]), .Z(n26) );
  CLKBUF_X1 U3 ( .A(SH[3]), .Z(n25) );
  CLKBUF_X1 U4 ( .A(SH[3]), .Z(n27) );
  CLKBUF_X1 U5 ( .A(SH[4]), .Z(n16) );
  CLKBUF_X1 U6 ( .A(SH[4]), .Z(n17) );
  CLKBUF_X1 U7 ( .A(SH[1]), .Z(n19) );
  CLKBUF_X1 U8 ( .A(SH[1]), .Z(n20) );
  CLKBUF_X1 U9 ( .A(SH[4]), .Z(n18) );
  CLKBUF_X1 U10 ( .A(SH[1]), .Z(n21) );
  CLKBUF_X1 U11 ( .A(SH[2]), .Z(n24) );
  CLKBUF_X1 U12 ( .A(SH[2]), .Z(n23) );
  CLKBUF_X1 U13 ( .A(SH[2]), .Z(n22) );
endmodule


module SHIFTER_GENERIC_N32_DW_lbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n18), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n18), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n18), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n18), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n18), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n18), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n18), .Z(B[25]) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n18), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n17), .Z(B[23]) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n17), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n17), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n17), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n17), .Z(B[19]) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n17), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n17), .Z(B[17]) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n17), .Z(B[16]) );
  MUX2_X1 M0_4_15 ( .A(\ML_int[4][15] ), .B(\ML_int[4][31] ), .S(n17), .Z(
        B[15]) );
  MUX2_X1 M0_4_14 ( .A(\ML_int[4][14] ), .B(\ML_int[4][30] ), .S(n17), .Z(
        B[14]) );
  MUX2_X1 M0_4_13 ( .A(\ML_int[4][13] ), .B(\ML_int[4][29] ), .S(n17), .Z(
        B[13]) );
  MUX2_X1 M0_4_12 ( .A(\ML_int[4][12] ), .B(\ML_int[4][28] ), .S(n17), .Z(
        B[12]) );
  MUX2_X1 M0_4_11 ( .A(\ML_int[4][11] ), .B(\ML_int[4][27] ), .S(n16), .Z(
        B[11]) );
  MUX2_X1 M0_4_10 ( .A(\ML_int[4][10] ), .B(\ML_int[4][26] ), .S(n16), .Z(
        B[10]) );
  MUX2_X1 M0_4_9 ( .A(\ML_int[4][9] ), .B(\ML_int[4][25] ), .S(n16), .Z(B[9])
         );
  MUX2_X1 M0_4_8 ( .A(\ML_int[4][8] ), .B(\ML_int[4][24] ), .S(n16), .Z(B[8])
         );
  MUX2_X1 M0_4_7 ( .A(\ML_int[4][7] ), .B(\ML_int[4][23] ), .S(n16), .Z(B[7])
         );
  MUX2_X1 M0_4_6 ( .A(\ML_int[4][6] ), .B(\ML_int[4][22] ), .S(n16), .Z(B[6])
         );
  MUX2_X1 M0_4_5 ( .A(\ML_int[4][5] ), .B(\ML_int[4][21] ), .S(n16), .Z(B[5])
         );
  MUX2_X1 M0_4_4 ( .A(\ML_int[4][4] ), .B(\ML_int[4][20] ), .S(n16), .Z(B[4])
         );
  MUX2_X1 M0_4_3 ( .A(\ML_int[4][3] ), .B(\ML_int[4][19] ), .S(n16), .Z(B[3])
         );
  MUX2_X1 M0_4_2 ( .A(\ML_int[4][2] ), .B(\ML_int[4][18] ), .S(n16), .Z(B[2])
         );
  MUX2_X1 M0_4_1 ( .A(\ML_int[4][1] ), .B(\ML_int[4][17] ), .S(n16), .Z(B[1])
         );
  MUX2_X1 M0_4_0 ( .A(\ML_int[4][0] ), .B(\ML_int[4][16] ), .S(n16), .Z(B[0])
         );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n27), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n27), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n27), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n27), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n27), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n27), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n27), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n27), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n26), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n26), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n26), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n26), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n26), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n26), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n26), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n26), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n26), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n26), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n26), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n26), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n25), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n25), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n25), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n25), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M0_3_7 ( .A(\ML_int[3][7] ), .B(\ML_int[3][31] ), .S(n25), .Z(
        \ML_int[4][7] ) );
  MUX2_X1 M0_3_6 ( .A(\ML_int[3][6] ), .B(\ML_int[3][30] ), .S(n25), .Z(
        \ML_int[4][6] ) );
  MUX2_X1 M0_3_5 ( .A(\ML_int[3][5] ), .B(\ML_int[3][29] ), .S(n25), .Z(
        \ML_int[4][5] ) );
  MUX2_X1 M0_3_4 ( .A(\ML_int[3][4] ), .B(\ML_int[3][28] ), .S(n25), .Z(
        \ML_int[4][4] ) );
  MUX2_X1 M0_3_3 ( .A(\ML_int[3][3] ), .B(\ML_int[3][27] ), .S(n25), .Z(
        \ML_int[4][3] ) );
  MUX2_X1 M0_3_2 ( .A(\ML_int[3][2] ), .B(\ML_int[3][26] ), .S(n25), .Z(
        \ML_int[4][2] ) );
  MUX2_X1 M0_3_1 ( .A(\ML_int[3][1] ), .B(\ML_int[3][25] ), .S(n25), .Z(
        \ML_int[4][1] ) );
  MUX2_X1 M0_3_0 ( .A(\ML_int[3][0] ), .B(\ML_int[3][24] ), .S(n25), .Z(
        \ML_int[4][0] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n24), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n24), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n24), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n24), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n24), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n24), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n24), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n24), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n22), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n22), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n22), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n22), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n22), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n22), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n22), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n22), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n22), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n22), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n22), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n22), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n23), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n23), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n23), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n23), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n23), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n23), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n23), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n23), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M0_2_3 ( .A(\ML_int[2][3] ), .B(\ML_int[2][31] ), .S(n23), .Z(
        \ML_int[3][3] ) );
  MUX2_X1 M0_2_2 ( .A(\ML_int[2][2] ), .B(\ML_int[2][30] ), .S(n23), .Z(
        \ML_int[3][2] ) );
  MUX2_X1 M0_2_1 ( .A(\ML_int[2][1] ), .B(\ML_int[2][29] ), .S(n23), .Z(
        \ML_int[3][1] ) );
  MUX2_X1 M0_2_0 ( .A(\ML_int[2][0] ), .B(\ML_int[2][28] ), .S(n23), .Z(
        \ML_int[3][0] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n21), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n21), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n21), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n21), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n21), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n21), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n21), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n21), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n19), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n19), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n19), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n19), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n19), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n19), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n19), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n19), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n19), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n19), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n19), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n19), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n20), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n20), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n20), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n20), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n20), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n20), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n20), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n20), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n20), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n20), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M0_1_1 ( .A(\ML_int[1][1] ), .B(\ML_int[1][31] ), .S(n20), .Z(
        \ML_int[2][1] ) );
  MUX2_X1 M0_1_0 ( .A(\ML_int[1][0] ), .B(\ML_int[1][30] ), .S(n20), .Z(
        \ML_int[2][0] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  MUX2_X1 M0_0_0 ( .A(A[0]), .B(A[31]), .S(SH[0]), .Z(\ML_int[1][0] ) );
  CLKBUF_X1 U2 ( .A(SH[3]), .Z(n25) );
  CLKBUF_X1 U3 ( .A(SH[3]), .Z(n26) );
  CLKBUF_X1 U4 ( .A(SH[3]), .Z(n27) );
  CLKBUF_X1 U5 ( .A(SH[4]), .Z(n16) );
  CLKBUF_X1 U6 ( .A(SH[4]), .Z(n17) );
  CLKBUF_X1 U7 ( .A(SH[1]), .Z(n19) );
  CLKBUF_X1 U8 ( .A(SH[1]), .Z(n20) );
  CLKBUF_X1 U9 ( .A(SH[4]), .Z(n18) );
  CLKBUF_X1 U10 ( .A(SH[1]), .Z(n21) );
  CLKBUF_X1 U11 ( .A(SH[2]), .Z(n24) );
  CLKBUF_X1 U12 ( .A(SH[2]), .Z(n23) );
  CLKBUF_X1 U13 ( .A(SH[2]), .Z(n22) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n45, n47, n48, n49, n50, n51, n52, n54, n56, n57, n58, n59, n60, n61,
         n63, n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n95, n96, n98, n99, n100, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n119,
         n122, n123, n125, n126, n129, n130, n131, n132, n133, n136, n138,
         n139, n140, n142, n144, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n172, n175, n176, n177, n182, n200,
         n202, n204, n208, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  MUX2_X1 U142 ( .A(\A[31] ), .B(A[30]), .S(n51), .Z(n84) );
  BUF_X2 U2 ( .A(n176), .Z(n182) );
  INV_X2 U3 ( .A(n182), .ZN(n177) );
  AOI221_X4 U4 ( .B1(n50), .B2(n213), .C1(n51), .C2(A[5]), .A(n96), .ZN(n32)
         );
  AOI221_X1 U5 ( .B1(n50), .B2(A[16]), .C1(n51), .C2(A[15]), .A(n140), .ZN(
        n109) );
  AOI221_X1 U6 ( .B1(n50), .B2(A[8]), .C1(n51), .C2(n211), .A(n52), .ZN(n20)
         );
  AOI221_X1 U7 ( .B1(n50), .B2(A[5]), .C1(n51), .C2(n220), .A(n169), .ZN(n35)
         );
  INV_X1 U8 ( .A(n38), .ZN(n6) );
  NAND2_X1 U9 ( .A1(n71), .A2(n177), .ZN(n38) );
  NAND2_X1 U10 ( .A1(n182), .A2(\A[31] ), .ZN(n58) );
  INV_X1 U11 ( .A(n3), .ZN(n41) );
  INV_X1 U12 ( .A(n100), .ZN(n74) );
  OAI21_X1 U13 ( .B1(n175), .B2(n69), .A(n58), .ZN(B[26]) );
  OAI21_X1 U14 ( .B1(n175), .B2(n67), .A(n58), .ZN(B[28]) );
  OAI21_X1 U15 ( .B1(n175), .B2(n68), .A(n58), .ZN(B[27]) );
  OAI21_X1 U16 ( .B1(n175), .B2(n14), .A(n58), .ZN(B[24]) );
  OAI21_X1 U17 ( .B1(n175), .B2(n21), .A(n58), .ZN(B[23]) );
  OAI21_X1 U18 ( .B1(n175), .B2(n59), .A(n58), .ZN(B[18]) );
  OAI21_X1 U19 ( .B1(n175), .B2(n107), .A(n58), .ZN(B[16]) );
  OAI21_X1 U20 ( .B1(n175), .B2(n90), .A(n58), .ZN(B[17]) );
  OAI21_X1 U21 ( .B1(n175), .B2(n4), .A(n58), .ZN(B[25]) );
  OAI21_X1 U22 ( .B1(n175), .B2(n66), .A(n58), .ZN(B[29]) );
  OAI21_X1 U23 ( .B1(n175), .B2(n57), .A(n58), .ZN(B[30]) );
  NOR2_X1 U24 ( .A1(n216), .A2(SH[3]), .ZN(n71) );
  INV_X1 U25 ( .A(n50), .ZN(n43) );
  INV_X1 U26 ( .A(n54), .ZN(n48) );
  INV_X1 U27 ( .A(n56), .ZN(n49) );
  INV_X1 U28 ( .A(n51), .ZN(n45) );
  NAND2_X1 U29 ( .A1(n73), .A2(n177), .ZN(n3) );
  AOI221_X1 U30 ( .B1(n75), .B2(n71), .C1(n76), .C2(n172), .A(n74), .ZN(n14)
         );
  AOI221_X1 U31 ( .B1(n84), .B2(n71), .C1(n79), .C2(n172), .A(n74), .ZN(n69)
         );
  AOI221_X1 U32 ( .B1(n77), .B2(n71), .C1(n78), .C2(n172), .A(n74), .ZN(n21)
         );
  AOI221_X1 U33 ( .B1(n70), .B2(n71), .C1(n72), .C2(n172), .A(n74), .ZN(n4) );
  AOI221_X1 U34 ( .B1(n80), .B2(n71), .C1(n31), .C2(n172), .A(n102), .ZN(n59)
         );
  INV_X1 U35 ( .A(n103), .ZN(n102) );
  AOI22_X1 U36 ( .A1(n104), .A2(n84), .B1(n83), .B2(n79), .ZN(n103) );
  AOI221_X1 U37 ( .B1(n11), .B2(n71), .C1(n9), .C2(n172), .A(n105), .ZN(n90)
         );
  INV_X1 U38 ( .A(n106), .ZN(n105) );
  AOI22_X1 U39 ( .A1(n104), .A2(n70), .B1(n83), .B2(n72), .ZN(n106) );
  AOI221_X1 U40 ( .B1(n18), .B2(n71), .C1(n17), .C2(n172), .A(n162), .ZN(n107)
         );
  INV_X1 U41 ( .A(n163), .ZN(n162) );
  AOI22_X1 U42 ( .A1(n104), .A2(n75), .B1(n83), .B2(n76), .ZN(n163) );
  AOI221_X1 U43 ( .B1(n76), .B2(n71), .C1(n18), .C2(n172), .A(n88), .ZN(n36)
         );
  INV_X1 U44 ( .A(n89), .ZN(n88) );
  AOI21_X1 U45 ( .B1(n83), .B2(n75), .A(n85), .ZN(n89) );
  AOI221_X1 U46 ( .B1(n79), .B2(n71), .C1(n80), .C2(n172), .A(n81), .ZN(n27)
         );
  INV_X1 U47 ( .A(n82), .ZN(n81) );
  AOI21_X1 U48 ( .B1(n83), .B2(n84), .A(n85), .ZN(n82) );
  AOI221_X1 U49 ( .B1(n72), .B2(n71), .C1(n11), .C2(n172), .A(n86), .ZN(n33)
         );
  INV_X1 U50 ( .A(n87), .ZN(n86) );
  AOI21_X1 U51 ( .B1(n83), .B2(n70), .A(n85), .ZN(n87) );
  AOI222_X1 U52 ( .A1(n6), .A2(n24), .B1(n8), .B2(n25), .C1(n10), .C2(n78), 
        .ZN(n133) );
  AOI222_X1 U53 ( .A1(n6), .A2(n17), .B1(n8), .B2(n18), .C1(n10), .C2(n76), 
        .ZN(n131) );
  OAI221_X1 U54 ( .B1(n26), .B2(n3), .C1(n27), .C2(n177), .A(n28), .ZN(B[6])
         );
  AOI222_X1 U55 ( .A1(n6), .A2(n29), .B1(n8), .B2(n30), .C1(n10), .C2(n31), 
        .ZN(n28) );
  OAI21_X1 U56 ( .B1(n175), .B2(n33), .A(n58), .ZN(B[21]) );
  OAI21_X1 U57 ( .B1(n175), .B2(n27), .A(n58), .ZN(B[22]) );
  OAI21_X1 U58 ( .B1(n175), .B2(n39), .A(n58), .ZN(B[19]) );
  OAI221_X1 U59 ( .B1(n43), .B2(n218), .C1(n45), .C2(n217), .A(n95), .ZN(n92)
         );
  NOR2_X1 U60 ( .A1(n100), .A2(n216), .ZN(n85) );
  BUF_X1 U61 ( .A(n73), .Z(n172) );
  AND2_X1 U62 ( .A1(n159), .A2(n216), .ZN(n8) );
  OAI221_X1 U63 ( .B1(n35), .B2(n3), .C1(n36), .C2(n177), .A(n37), .ZN(B[4])
         );
  AOI222_X1 U64 ( .A1(n6), .A2(n19), .B1(n8), .B2(n16), .C1(n10), .C2(n17), 
        .ZN(n37) );
  OAI221_X1 U65 ( .B1(n20), .B2(n3), .C1(n21), .C2(n177), .A(n22), .ZN(B[7])
         );
  AOI222_X1 U66 ( .A1(n6), .A2(n23), .B1(n8), .B2(n24), .C1(n10), .C2(n25), 
        .ZN(n22) );
  OAI221_X1 U67 ( .B1(n13), .B2(n3), .C1(n14), .C2(n177), .A(n15), .ZN(B[8])
         );
  INV_X1 U68 ( .A(n19), .ZN(n13) );
  AOI222_X1 U69 ( .A1(n6), .A2(n16), .B1(n8), .B2(n17), .C1(n10), .C2(n18), 
        .ZN(n15) );
  OAI221_X1 U70 ( .B1(n32), .B2(n3), .C1(n33), .C2(n177), .A(n34), .ZN(B[5])
         );
  AOI222_X1 U71 ( .A1(n6), .A2(n12), .B1(n8), .B2(n7), .C1(n10), .C2(n9), .ZN(
        n34) );
  OAI221_X1 U72 ( .B1(n2), .B2(n3), .C1(n4), .C2(n177), .A(n5), .ZN(B[9]) );
  INV_X1 U73 ( .A(n12), .ZN(n2) );
  AOI222_X1 U74 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .C1(n10), .C2(n11), .ZN(
        n5) );
  OAI221_X1 U75 ( .B1(n148), .B2(n3), .C1(n69), .C2(n177), .A(n149), .ZN(B[10]) );
  INV_X1 U76 ( .A(n29), .ZN(n148) );
  AOI222_X1 U77 ( .A1(n6), .A2(n30), .B1(n8), .B2(n31), .C1(n10), .C2(n80), 
        .ZN(n149) );
  OAI221_X1 U78 ( .B1(n115), .B2(n3), .C1(n66), .C2(n177), .A(n116), .ZN(B[13]) );
  INV_X1 U79 ( .A(n7), .ZN(n115) );
  AOI222_X1 U80 ( .A1(n6), .A2(n9), .B1(n8), .B2(n11), .C1(n10), .C2(n72), 
        .ZN(n116) );
  OAI221_X1 U81 ( .B1(n32), .B2(n38), .C1(n90), .C2(n177), .A(n91), .ZN(B[1])
         );
  AOI222_X1 U82 ( .A1(n10), .A2(n7), .B1(n41), .B2(n92), .C1(n8), .C2(n12), 
        .ZN(n91) );
  OAI221_X1 U83 ( .B1(n108), .B2(n38), .C1(n109), .C2(n3), .A(n110), .ZN(B[15]) );
  INV_X1 U84 ( .A(n25), .ZN(n108) );
  AOI221_X1 U85 ( .B1(n10), .B2(n77), .C1(n8), .C2(n78), .A(n111), .ZN(n110)
         );
  INV_X1 U86 ( .A(n58), .ZN(n111) );
  AND2_X1 U87 ( .A1(SH[3]), .A2(n216), .ZN(n83) );
  AOI21_X1 U88 ( .B1(n77), .B2(n172), .A(n114), .ZN(n68) );
  AOI21_X1 U89 ( .B1(n75), .B2(n172), .A(n114), .ZN(n67) );
  NAND2_X1 U90 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n100) );
  AOI221_X1 U91 ( .B1(n78), .B2(n71), .C1(n25), .C2(n172), .A(n98), .ZN(n39)
         );
  INV_X1 U92 ( .A(n99), .ZN(n98) );
  AOI21_X1 U93 ( .B1(n83), .B2(n77), .A(n85), .ZN(n99) );
  INV_X1 U94 ( .A(n112), .ZN(n30) );
  INV_X1 U95 ( .A(n109), .ZN(n24) );
  OAI21_X1 U96 ( .B1(n175), .B2(n36), .A(n58), .ZN(B[20]) );
  OAI221_X1 U97 ( .B1(n26), .B2(n38), .C1(n59), .C2(n177), .A(n60), .ZN(B[2])
         );
  AOI222_X1 U98 ( .A1(n10), .A2(n30), .B1(n41), .B2(n61), .C1(n8), .C2(n29), 
        .ZN(n60) );
  OAI221_X1 U99 ( .B1(n132), .B2(n3), .C1(n68), .C2(n177), .A(n133), .ZN(B[11]) );
  INV_X1 U100 ( .A(n23), .ZN(n132) );
  OAI221_X1 U101 ( .B1(n130), .B2(n3), .C1(n67), .C2(n177), .A(n131), .ZN(
        B[12]) );
  INV_X1 U102 ( .A(n16), .ZN(n130) );
  OAI221_X1 U103 ( .B1(n35), .B2(n38), .C1(n107), .C2(n177), .A(n156), .ZN(
        B[0]) );
  AOI222_X1 U104 ( .A1(n10), .A2(n16), .B1(n41), .B2(n157), .C1(n8), .C2(n19), 
        .ZN(n156) );
  AND2_X1 U105 ( .A1(SH[3]), .A2(n177), .ZN(n159) );
  OAI221_X1 U106 ( .B1(n112), .B2(n3), .C1(n57), .C2(n177), .A(n113), .ZN(
        B[14]) );
  AOI222_X1 U107 ( .A1(n6), .A2(n31), .B1(n8), .B2(n80), .C1(n10), .C2(n79), 
        .ZN(n113) );
  AOI221_X1 U108 ( .B1(n50), .B2(n211), .C1(n51), .C2(n213), .A(n64), .ZN(n26)
         );
  OAI22_X1 U109 ( .A1(n222), .A2(n54), .B1(n223), .B2(n56), .ZN(n64) );
  OAI21_X1 U110 ( .B1(n216), .B2(n210), .A(n100), .ZN(n114) );
  AOI21_X1 U111 ( .B1(n70), .B2(n172), .A(n114), .ZN(n66) );
  AOI21_X1 U112 ( .B1(n84), .B2(n172), .A(n114), .ZN(n57) );
  OAI221_X1 U113 ( .B1(n43), .B2(n165), .C1(n45), .C2(n142), .A(n166), .ZN(n75) );
  INV_X1 U114 ( .A(A[29]), .ZN(n165) );
  AOI22_X1 U115 ( .A1(A[30]), .A2(n48), .B1(\A[31] ), .B2(n49), .ZN(n166) );
  OAI221_X1 U116 ( .B1(n43), .B2(n232), .C1(n45), .C2(n204), .A(n136), .ZN(n78) );
  AOI22_X1 U117 ( .A1(A[25]), .A2(n48), .B1(A[26]), .B2(n49), .ZN(n136) );
  OAI221_X1 U118 ( .B1(n43), .B2(n208), .C1(n45), .C2(n234), .A(n154), .ZN(n79) );
  AOI22_X1 U119 ( .A1(A[28]), .A2(n48), .B1(A[29]), .B2(n49), .ZN(n154) );
  OAI221_X1 U120 ( .B1(n43), .B2(n234), .C1(n45), .C2(n233), .A(n119), .ZN(n72) );
  AOI22_X1 U121 ( .A1(A[27]), .A2(n48), .B1(A[28]), .B2(n49), .ZN(n119) );
  OAI221_X1 U122 ( .B1(n43), .B2(n233), .C1(n45), .C2(n232), .A(n164), .ZN(n76) );
  AOI22_X1 U123 ( .A1(A[26]), .A2(n48), .B1(A[27]), .B2(n49), .ZN(n164) );
  OAI221_X1 U124 ( .B1(n43), .B2(n204), .C1(n45), .C2(n231), .A(n150), .ZN(n80) );
  AOI22_X1 U125 ( .A1(A[24]), .A2(n48), .B1(A[25]), .B2(n49), .ZN(n150) );
  OAI221_X1 U126 ( .B1(n43), .B2(n231), .C1(n45), .C2(n202), .A(n122), .ZN(n11) );
  AOI22_X1 U127 ( .A1(A[23]), .A2(n48), .B1(A[24]), .B2(n49), .ZN(n122) );
  OAI221_X1 U128 ( .B1(n43), .B2(n202), .C1(n230), .C2(n45), .A(n168), .ZN(n18) );
  AOI22_X1 U129 ( .A1(A[22]), .A2(n48), .B1(A[23]), .B2(n49), .ZN(n168) );
  OAI221_X1 U130 ( .B1(n43), .B2(n229), .C1(n45), .C2(n227), .A(n129), .ZN(n7)
         );
  AOI22_X1 U131 ( .A1(A[15]), .A2(n48), .B1(A[16]), .B2(n49), .ZN(n129) );
  OAI221_X1 U132 ( .B1(n43), .B2(n227), .C1(n45), .C2(n226), .A(n161), .ZN(n16) );
  AOI22_X1 U133 ( .A1(n228), .A2(n48), .B1(A[15]), .B2(n49), .ZN(n161) );
  OAI221_X1 U134 ( .B1(n43), .B2(n123), .C1(n45), .C2(n200), .A(n125), .ZN(n9)
         );
  AOI22_X1 U135 ( .A1(A[19]), .A2(n48), .B1(A[20]), .B2(n49), .ZN(n125) );
  OAI221_X1 U136 ( .B1(n43), .B2(n142), .C1(n45), .C2(n208), .A(n144), .ZN(n77) );
  AOI22_X1 U137 ( .A1(A[29]), .A2(n48), .B1(A[30]), .B2(n49), .ZN(n144) );
  OAI221_X1 U138 ( .B1(n230), .B2(n43), .C1(n138), .C2(n45), .A(n139), .ZN(n25) );
  AOI22_X1 U139 ( .A1(A[21]), .A2(n48), .B1(A[22]), .B2(n49), .ZN(n139) );
  OAI221_X1 U140 ( .B1(n54), .B2(n123), .C1(n138), .C2(n56), .A(n167), .ZN(n17) );
  AOI22_X1 U141 ( .A1(A[17]), .A2(n50), .B1(A[16]), .B2(n51), .ZN(n167) );
  OAI221_X1 U143 ( .B1(n138), .B2(n43), .C1(n123), .C2(n45), .A(n151), .ZN(n31) );
  AOI22_X1 U144 ( .A1(A[20]), .A2(n48), .B1(A[21]), .B2(n49), .ZN(n151) );
  OAI221_X1 U145 ( .B1(n43), .B2(n225), .C1(n45), .C2(n224), .A(n155), .ZN(n29) );
  AOI22_X1 U146 ( .A1(A[12]), .A2(n48), .B1(A[13]), .B2(n49), .ZN(n155) );
  OAI221_X1 U147 ( .B1(n43), .B2(n224), .C1(n45), .C2(n223), .A(n93), .ZN(n12)
         );
  AOI22_X1 U148 ( .A1(A[11]), .A2(n48), .B1(A[12]), .B2(n49), .ZN(n93) );
  OAI221_X1 U149 ( .B1(n43), .B2(n226), .C1(n45), .C2(n225), .A(n147), .ZN(n23) );
  AOI22_X1 U150 ( .A1(A[13]), .A2(n48), .B1(n228), .B2(n49), .ZN(n147) );
  AOI221_X1 U151 ( .B1(n50), .B2(A[15]), .C1(n51), .C2(n228), .A(n152), .ZN(
        n112) );
  INV_X1 U152 ( .A(n153), .ZN(n152) );
  AOI22_X1 U153 ( .A1(A[16]), .A2(n48), .B1(A[17]), .B2(n49), .ZN(n153) );
  OAI22_X1 U154 ( .A1(n200), .A2(n54), .B1(n123), .B2(n56), .ZN(n140) );
  OAI221_X1 U155 ( .B1(n43), .B2(n219), .C1(n45), .C2(n218), .A(n63), .ZN(n61)
         );
  OAI221_X1 U156 ( .B1(n20), .B2(n38), .C1(n39), .C2(n177), .A(n40), .ZN(B[3])
         );
  AOI222_X1 U157 ( .A1(n10), .A2(n24), .B1(n41), .B2(n42), .C1(n8), .C2(n23), 
        .ZN(n40) );
  OAI221_X1 U158 ( .B1(n43), .B2(n221), .C1(n45), .C2(n219), .A(n47), .ZN(n42)
         );
  OAI221_X1 U159 ( .B1(n43), .B2(n223), .C1(n45), .C2(n222), .A(n158), .ZN(n19) );
  AOI22_X1 U160 ( .A1(A[10]), .A2(n48), .B1(A[11]), .B2(n49), .ZN(n158) );
  INV_X1 U161 ( .A(A[18]), .ZN(n123) );
  INV_X1 U162 ( .A(n126), .ZN(n70) );
  INV_X1 U163 ( .A(A[19]), .ZN(n138) );
  INV_X1 U164 ( .A(A[23]), .ZN(n204) );
  INV_X1 U165 ( .A(A[21]), .ZN(n202) );
  INV_X1 U166 ( .A(A[28]), .ZN(n142) );
  INV_X1 U167 ( .A(A[17]), .ZN(n200) );
  INV_X1 U168 ( .A(A[27]), .ZN(n208) );
  INV_X1 U169 ( .A(\A[31] ), .ZN(n210) );
  CLKBUF_X1 U170 ( .A(SH[4]), .Z(n176) );
  OAI221_X1 U171 ( .B1(n54), .B2(n218), .C1(n56), .C2(n219), .A(n160), .ZN(
        n157) );
  OAI22_X1 U172 ( .A1(n212), .A2(n54), .B1(n222), .B2(n56), .ZN(n96) );
  OAI22_X1 U173 ( .A1(n214), .A2(n54), .B1(n212), .B2(n56), .ZN(n169) );
  OAI22_X1 U174 ( .A1(n223), .A2(n54), .B1(n224), .B2(n56), .ZN(n52) );
  CLKBUF_X1 U175 ( .A(SH[4]), .Z(n175) );
  AOI22_X1 U176 ( .A1(A[1]), .A2(n50), .B1(A[0]), .B2(n51), .ZN(n160) );
  AOI22_X1 U177 ( .A1(A[3]), .A2(n48), .B1(n220), .B2(n49), .ZN(n95) );
  AOI22_X1 U178 ( .A1(A[5]), .A2(n48), .B1(n213), .B2(n49), .ZN(n47) );
  AOI22_X1 U179 ( .A1(n220), .A2(n48), .B1(A[5]), .B2(n49), .ZN(n63) );
  INV_X1 U180 ( .A(A[7]), .ZN(n212) );
  AND2_X1 U181 ( .A1(SH[2]), .A2(SH[3]), .ZN(n104) );
  AOI222_X1 U182 ( .A1(n51), .A2(A[29]), .B1(n50), .B2(A[30]), .C1(SH[1]), 
        .C2(\A[31] ), .ZN(n126) );
  NOR2_X1 U183 ( .A1(SH[0]), .A2(SH[1]), .ZN(n51) );
  NOR2_X1 U184 ( .A1(n215), .A2(SH[1]), .ZN(n50) );
  NAND2_X1 U185 ( .A1(SH[1]), .A2(n215), .ZN(n54) );
  NAND2_X1 U186 ( .A1(SH[0]), .A2(SH[1]), .ZN(n56) );
  AND2_X1 U187 ( .A1(SH[2]), .A2(n159), .ZN(n10) );
  NOR2_X1 U188 ( .A1(SH[2]), .A2(SH[3]), .ZN(n73) );
  INV_X1 U189 ( .A(n212), .ZN(n211) );
  INV_X1 U190 ( .A(n214), .ZN(n213) );
  INV_X1 U191 ( .A(A[6]), .ZN(n214) );
  INV_X1 U192 ( .A(SH[0]), .ZN(n215) );
  INV_X1 U193 ( .A(SH[2]), .ZN(n216) );
  INV_X1 U194 ( .A(A[1]), .ZN(n217) );
  INV_X1 U195 ( .A(A[2]), .ZN(n218) );
  INV_X1 U196 ( .A(A[3]), .ZN(n219) );
  INV_X1 U197 ( .A(n221), .ZN(n220) );
  INV_X1 U198 ( .A(A[4]), .ZN(n221) );
  INV_X1 U199 ( .A(A[8]), .ZN(n222) );
  INV_X1 U200 ( .A(A[9]), .ZN(n223) );
  INV_X1 U201 ( .A(A[10]), .ZN(n224) );
  INV_X1 U202 ( .A(A[11]), .ZN(n225) );
  INV_X1 U203 ( .A(A[12]), .ZN(n226) );
  INV_X1 U204 ( .A(A[13]), .ZN(n227) );
  INV_X1 U205 ( .A(n229), .ZN(n228) );
  INV_X1 U206 ( .A(A[14]), .ZN(n229) );
  INV_X1 U207 ( .A(A[20]), .ZN(n230) );
  INV_X1 U208 ( .A(A[22]), .ZN(n231) );
  INV_X1 U209 ( .A(A[24]), .ZN(n232) );
  INV_X1 U210 ( .A(A[25]), .ZN(n233) );
  INV_X1 U211 ( .A(A[26]), .ZN(n234) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n48, n50, n51, n52, n53, n54, n55, n57, n59, n60, n61, n62, n63, n64,
         n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n110,
         n111, n113, n114, n116, n118, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n132, n133, n136, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n151, n153, n155, n156,
         n157, n158, n159, n161, n162, n164, n165, n166, n167, n168, n174,
         n175, n176, n177, n178, n180, n202, n203, n205, n206, n207, n208,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240;

  MUX2_X1 U104 ( .A(n77), .B(n60), .S(SH[2]), .Z(n91) );
  BUF_X2 U3 ( .A(n178), .Z(n176) );
  BUF_X2 U4 ( .A(n178), .Z(n177) );
  INV_X2 U5 ( .A(n177), .ZN(n180) );
  AOI221_X1 U6 ( .B1(n53), .B2(A[7]), .C1(n54), .C2(A[6]), .A(n162), .ZN(n36)
         );
  NOR2_X1 U7 ( .A1(n218), .A2(SH[3]), .ZN(n75) );
  INV_X1 U8 ( .A(n5), .ZN(n43) );
  NAND2_X1 U9 ( .A1(n74), .A2(n180), .ZN(n5) );
  INV_X1 U10 ( .A(n40), .ZN(n8) );
  INV_X1 U11 ( .A(n167), .ZN(n54) );
  NAND2_X1 U12 ( .A1(n75), .A2(n180), .ZN(n40) );
  NOR2_X1 U13 ( .A1(n180), .A2(n125), .ZN(n101) );
  INV_X1 U14 ( .A(n125), .ZN(n74) );
  NOR3_X1 U15 ( .A1(n71), .A2(n174), .A3(SH[3]), .ZN(B[27]) );
  NOR2_X1 U16 ( .A1(n219), .A2(n174), .ZN(n148) );
  NOR2_X1 U17 ( .A1(n174), .A2(n72), .ZN(B[26]) );
  INV_X1 U18 ( .A(n4), .ZN(n35) );
  INV_X1 U19 ( .A(n14), .ZN(n39) );
  NOR2_X1 U20 ( .A1(n175), .A2(n82), .ZN(B[17]) );
  NOR2_X1 U21 ( .A1(n177), .A2(n62), .ZN(B[18]) );
  NOR2_X1 U22 ( .A1(n174), .A2(n97), .ZN(B[16]) );
  NOR2_X1 U23 ( .A1(n175), .A2(n21), .ZN(B[23]) );
  NOR2_X1 U24 ( .A1(n176), .A2(n41), .ZN(B[19]) );
  NOR2_X1 U25 ( .A1(n176), .A2(n33), .ZN(B[21]) );
  NOR2_X1 U26 ( .A1(n176), .A2(n27), .ZN(B[22]) );
  NOR2_X1 U27 ( .A1(n176), .A2(n37), .ZN(B[20]) );
  NOR2_X1 U28 ( .A1(n175), .A2(n6), .ZN(B[25]) );
  AND2_X1 U29 ( .A1(n69), .A2(n43), .ZN(B[29]) );
  INV_X1 U30 ( .A(n122), .ZN(B[12]) );
  OAI221_X1 U31 ( .B1(n20), .B2(n5), .C1(n21), .C2(n180), .A(n22), .ZN(B[7])
         );
  OAI221_X1 U32 ( .B1(n14), .B2(n5), .C1(n15), .C2(n180), .A(n16), .ZN(B[8])
         );
  AND2_X1 U33 ( .A1(n61), .A2(n43), .ZN(B[30]) );
  AND2_X1 U34 ( .A1(n43), .A2(n60), .ZN(B[31]) );
  NOR2_X1 U35 ( .A1(n175), .A2(n15), .ZN(B[24]) );
  OAI222_X1 U36 ( .A1(n57), .A2(n111), .B1(n168), .B2(n213), .C1(n59), .C2(
        n113), .ZN(n69) );
  INV_X1 U37 ( .A(n46), .ZN(n53) );
  INV_X1 U38 ( .A(n52), .ZN(n59) );
  OAI22_X1 U39 ( .A1(n59), .A2(n111), .B1(n57), .B2(n213), .ZN(n61) );
  AOI222_X1 U40 ( .A1(n73), .A2(n75), .B1(n69), .B2(n78), .C1(n13), .C2(n74), 
        .ZN(n33) );
  AOI222_X1 U41 ( .A1(n77), .A2(n75), .B1(n60), .B2(n78), .C1(n79), .C2(n74), 
        .ZN(n21) );
  AOI222_X1 U42 ( .A1(n80), .A2(n75), .B1(n61), .B2(n78), .C1(n81), .C2(n74), 
        .ZN(n27) );
  AOI222_X1 U43 ( .A1(n76), .A2(n75), .B1(n70), .B2(n78), .C1(n19), .C2(n74), 
        .ZN(n37) );
  AOI222_X1 U44 ( .A1(n25), .A2(n74), .B1(n79), .B2(n75), .C1(n91), .C2(SH[3]), 
        .ZN(n41) );
  INV_X1 U45 ( .A(n51), .ZN(n57) );
  AOI221_X1 U46 ( .B1(n53), .B2(n227), .C1(n54), .C2(n225), .A(n68), .ZN(n26)
         );
  OAI22_X1 U47 ( .A1(n214), .A2(n57), .B1(n215), .B2(n59), .ZN(n68) );
  AOI221_X1 U48 ( .B1(n53), .B2(n229), .C1(n54), .C2(n227), .A(n55), .ZN(n20)
         );
  OAI22_X1 U49 ( .A1(n226), .A2(n57), .B1(n214), .B2(n59), .ZN(n55) );
  AOI221_X1 U50 ( .B1(n53), .B2(n233), .C1(n54), .C2(n231), .A(n85), .ZN(n4)
         );
  OAI22_X1 U51 ( .A1(n230), .A2(n57), .B1(n228), .B2(n59), .ZN(n85) );
  AOI221_X1 U52 ( .B1(n53), .B2(n231), .C1(n54), .C2(n229), .A(n147), .ZN(n14)
         );
  OAI22_X1 U53 ( .A1(n228), .A2(n57), .B1(n226), .B2(n59), .ZN(n147) );
  AOI221_X1 U54 ( .B1(n19), .B2(n75), .C1(n18), .C2(n74), .A(n155), .ZN(n97)
         );
  INV_X1 U55 ( .A(n156), .ZN(n155) );
  AOI22_X1 U56 ( .A1(n94), .A2(n70), .B1(n78), .B2(n76), .ZN(n156) );
  AOI221_X1 U57 ( .B1(n81), .B2(n75), .C1(n31), .C2(n74), .A(n92), .ZN(n62) );
  INV_X1 U58 ( .A(n93), .ZN(n92) );
  AOI22_X1 U59 ( .A1(n94), .A2(n61), .B1(n78), .B2(n80), .ZN(n93) );
  AOI222_X1 U60 ( .A1(n8), .A2(n17), .B1(n10), .B2(n18), .C1(n12), .C2(n19), 
        .ZN(n16) );
  AOI222_X1 U61 ( .A1(n12), .A2(n73), .B1(n101), .B2(n69), .C1(n10), .C2(n13), 
        .ZN(n107) );
  AOI222_X1 U62 ( .A1(n12), .A2(n80), .B1(n101), .B2(n61), .C1(n10), .C2(n81), 
        .ZN(n104) );
  AOI222_X1 U63 ( .A1(n12), .A2(n77), .B1(n101), .B2(n60), .C1(n10), .C2(n79), 
        .ZN(n100) );
  AOI222_X1 U64 ( .A1(n8), .A2(n23), .B1(n10), .B2(n24), .C1(n12), .C2(n25), 
        .ZN(n22) );
  AOI221_X1 U65 ( .B1(n12), .B2(n79), .C1(n10), .C2(n25), .A(n127), .ZN(n126)
         );
  NOR3_X1 U66 ( .A1(n180), .A2(SH[3]), .A3(n71), .ZN(n127) );
  AOI221_X1 U67 ( .B1(n18), .B2(n8), .C1(n17), .C2(n43), .A(n123), .ZN(n122)
         );
  INV_X1 U68 ( .A(n124), .ZN(n123) );
  AOI222_X1 U69 ( .A1(n12), .A2(n76), .B1(n101), .B2(n70), .C1(n10), .C2(n19), 
        .ZN(n124) );
  BUF_X1 U70 ( .A(n52), .Z(n164) );
  INV_X1 U71 ( .A(n165), .ZN(n166) );
  INV_X1 U72 ( .A(n51), .ZN(n165) );
  AND2_X1 U73 ( .A1(n148), .A2(n218), .ZN(n10) );
  OAI221_X1 U74 ( .B1(n65), .B2(n5), .C1(n72), .C2(n180), .A(n139), .ZN(B[10])
         );
  AOI222_X1 U75 ( .A1(n8), .A2(n30), .B1(n10), .B2(n31), .C1(n12), .C2(n81), 
        .ZN(n139) );
  OAI221_X1 U76 ( .B1(n36), .B2(n5), .C1(n37), .C2(n180), .A(n38), .ZN(B[4])
         );
  AOI222_X1 U77 ( .A1(n8), .A2(n39), .B1(n10), .B2(n17), .C1(n12), .C2(n18), 
        .ZN(n38) );
  OAI221_X1 U78 ( .B1(n32), .B2(n5), .C1(n33), .C2(n180), .A(n34), .ZN(B[5])
         );
  AOI222_X1 U79 ( .A1(n8), .A2(n35), .B1(n10), .B2(n9), .C1(n12), .C2(n11), 
        .ZN(n34) );
  OAI221_X1 U80 ( .B1(n26), .B2(n5), .C1(n27), .C2(n180), .A(n28), .ZN(B[6])
         );
  AOI222_X1 U81 ( .A1(n8), .A2(n29), .B1(n10), .B2(n30), .C1(n12), .C2(n31), 
        .ZN(n28) );
  AOI22_X1 U82 ( .A1(n80), .A2(n74), .B1(n61), .B2(n75), .ZN(n72) );
  AOI22_X1 U83 ( .A1(n76), .A2(n74), .B1(n70), .B2(n75), .ZN(n15) );
  AOI22_X1 U84 ( .A1(n73), .A2(n74), .B1(n69), .B2(n75), .ZN(n6) );
  OAI221_X1 U85 ( .B1(n4), .B2(n5), .C1(n6), .C2(n180), .A(n7), .ZN(B[9]) );
  AOI222_X1 U86 ( .A1(n8), .A2(n9), .B1(n10), .B2(n11), .C1(n12), .C2(n13), 
        .ZN(n7) );
  NOR2_X1 U87 ( .A1(n213), .A2(n59), .ZN(n60) );
  OAI221_X1 U88 ( .B1(n26), .B2(n40), .C1(n62), .C2(n180), .A(n63), .ZN(B[2])
         );
  AOI222_X1 U89 ( .A1(n12), .A2(n30), .B1(n43), .B2(n64), .C1(n10), .C2(n29), 
        .ZN(n63) );
  OAI221_X1 U90 ( .B1(n46), .B2(n224), .C1(n168), .C2(n223), .A(n67), .ZN(n64)
         );
  OAI221_X1 U91 ( .B1(n32), .B2(n40), .C1(n82), .C2(n180), .A(n83), .ZN(B[1])
         );
  AOI222_X1 U92 ( .A1(n12), .A2(n9), .B1(n43), .B2(n84), .C1(n10), .C2(n35), 
        .ZN(n83) );
  OAI221_X1 U93 ( .B1(n46), .B2(n223), .C1(n168), .C2(n222), .A(n89), .ZN(n84)
         );
  NOR2_X1 U94 ( .A1(n218), .A2(n219), .ZN(n94) );
  BUF_X1 U95 ( .A(n48), .Z(n167) );
  BUF_X1 U96 ( .A(n48), .Z(n168) );
  INV_X1 U97 ( .A(SH[3]), .ZN(n219) );
  BUF_X1 U98 ( .A(n176), .Z(n174) );
  NAND2_X1 U99 ( .A1(n218), .A2(n219), .ZN(n125) );
  INV_X1 U100 ( .A(n24), .ZN(n99) );
  INV_X1 U101 ( .A(n11), .ZN(n105) );
  INV_X1 U102 ( .A(n208), .ZN(n207) );
  INV_X1 U103 ( .A(n206), .ZN(n205) );
  INV_X1 U105 ( .A(n65), .ZN(n29) );
  INV_X1 U106 ( .A(n45), .ZN(n23) );
  INV_X1 U107 ( .A(n31), .ZN(n102) );
  AOI221_X1 U108 ( .B1(n13), .B2(n75), .C1(n11), .C2(n74), .A(n95), .ZN(n82)
         );
  INV_X1 U109 ( .A(n96), .ZN(n95) );
  AOI22_X1 U110 ( .A1(n94), .A2(n69), .B1(n78), .B2(n73), .ZN(n96) );
  INV_X1 U111 ( .A(n91), .ZN(n71) );
  AND2_X1 U112 ( .A1(n70), .A2(n43), .ZN(B[28]) );
  OAI221_X1 U113 ( .B1(n36), .B2(n40), .C1(n97), .C2(n180), .A(n145), .ZN(B[0]) );
  OAI221_X1 U114 ( .B1(n99), .B2(n40), .C1(n45), .C2(n5), .A(n126), .ZN(B[11])
         );
  OAI221_X1 U115 ( .B1(n105), .B2(n40), .C1(n106), .C2(n5), .A(n107), .ZN(
        B[13]) );
  INV_X1 U116 ( .A(n9), .ZN(n106) );
  OAI221_X1 U117 ( .B1(n98), .B2(n40), .C1(n99), .C2(n5), .A(n100), .ZN(B[15])
         );
  INV_X1 U118 ( .A(n25), .ZN(n98) );
  OAI221_X1 U119 ( .B1(n102), .B2(n40), .C1(n103), .C2(n5), .A(n104), .ZN(
        B[14]) );
  INV_X1 U120 ( .A(n30), .ZN(n103) );
  CLKBUF_X1 U121 ( .A(n176), .Z(n175) );
  OAI22_X1 U122 ( .A1(n224), .A2(n57), .B1(n223), .B2(n59), .ZN(n162) );
  OAI221_X1 U123 ( .B1(n46), .B2(n213), .C1(n167), .C2(n111), .A(n158), .ZN(
        n70) );
  AOI22_X1 U124 ( .A1(A[29]), .A2(n166), .B1(A[28]), .B2(n164), .ZN(n158) );
  OAI221_X1 U125 ( .B1(n46), .B2(n237), .C1(n167), .C2(n120), .A(n121), .ZN(
        n11) );
  AOI22_X1 U126 ( .A1(A[18]), .A2(n166), .B1(A[17]), .B2(n164), .ZN(n121) );
  OAI221_X1 U127 ( .B1(n46), .B2(n120), .C1(n167), .C2(n136), .A(n159), .ZN(
        n18) );
  AOI22_X1 U128 ( .A1(A[17]), .A2(n166), .B1(A[16]), .B2(n164), .ZN(n159) );
  OAI221_X1 U129 ( .B1(n46), .B2(n203), .C1(n168), .C2(n202), .A(n142), .ZN(
        n30) );
  AOI22_X1 U130 ( .A1(A[15]), .A2(n166), .B1(n235), .B2(n164), .ZN(n142) );
  OAI221_X1 U131 ( .B1(n46), .B2(n202), .C1(n168), .C2(n216), .A(n118), .ZN(n9) );
  AOI22_X1 U132 ( .A1(n235), .A2(n166), .B1(A[13]), .B2(n164), .ZN(n118) );
  OAI221_X1 U133 ( .B1(n46), .B2(n216), .C1(n168), .C2(n236), .A(n153), .ZN(
        n17) );
  AOI22_X1 U134 ( .A1(A[13]), .A2(n166), .B1(n233), .B2(n164), .ZN(n153) );
  OAI221_X1 U135 ( .B1(n46), .B2(n114), .C1(n168), .C2(n212), .A(n116), .ZN(
        n73) );
  AOI22_X1 U136 ( .A1(A[26]), .A2(n166), .B1(A[25]), .B2(n164), .ZN(n116) );
  OAI221_X1 U137 ( .B1(n46), .B2(n212), .C1(n167), .C2(n240), .A(n157), .ZN(
        n76) );
  AOI22_X1 U138 ( .A1(A[25]), .A2(n166), .B1(A[24]), .B2(n164), .ZN(n157) );
  OAI221_X1 U139 ( .B1(n46), .B2(n113), .C1(n168), .C2(n114), .A(n143), .ZN(
        n80) );
  AOI22_X1 U140 ( .A1(A[27]), .A2(n166), .B1(A[26]), .B2(n164), .ZN(n143) );
  OAI221_X1 U141 ( .B1(n46), .B2(n239), .C1(n168), .C2(n238), .A(n140), .ZN(
        n81) );
  AOI22_X1 U142 ( .A1(n207), .A2(n166), .B1(A[22]), .B2(n164), .ZN(n140) );
  OAI221_X1 U143 ( .B1(n46), .B2(n238), .C1(n168), .C2(n208), .A(n110), .ZN(
        n13) );
  AOI22_X1 U144 ( .A1(A[22]), .A2(n166), .B1(n205), .B2(n164), .ZN(n110) );
  OAI221_X1 U145 ( .B1(n46), .B2(n240), .C1(n167), .C2(n239), .A(n132), .ZN(
        n79) );
  AOI22_X1 U146 ( .A1(A[24]), .A2(n166), .B1(n207), .B2(n164), .ZN(n132) );
  OAI221_X1 U147 ( .B1(n46), .B2(n136), .C1(n168), .C2(n203), .A(n138), .ZN(
        n24) );
  AOI22_X1 U148 ( .A1(A[16]), .A2(n166), .B1(A[15]), .B2(n164), .ZN(n138) );
  OAI221_X1 U149 ( .B1(n46), .B2(n111), .C1(n167), .C2(n113), .A(n128), .ZN(
        n77) );
  AOI22_X1 U150 ( .A1(A[28]), .A2(n51), .B1(A[27]), .B2(n52), .ZN(n128) );
  OAI221_X1 U151 ( .B1(n237), .B2(n57), .C1(n120), .C2(n59), .A(n129), .ZN(n25) );
  AOI22_X1 U152 ( .A1(A[22]), .A2(n53), .B1(n205), .B2(n54), .ZN(n129) );
  OAI221_X1 U153 ( .B1(n120), .B2(n57), .C1(n136), .C2(n59), .A(n141), .ZN(n31) );
  AOI22_X1 U154 ( .A1(n205), .A2(n53), .B1(n54), .B2(A[20]), .ZN(n141) );
  OAI221_X1 U155 ( .B1(n57), .B2(n206), .C1(n237), .C2(n59), .A(n161), .ZN(n19) );
  AOI22_X1 U156 ( .A1(n207), .A2(n53), .B1(A[22]), .B2(n54), .ZN(n161) );
  AOI221_X1 U157 ( .B1(n53), .B2(A[13]), .C1(n54), .C2(n233), .A(n144), .ZN(
        n65) );
  OAI22_X1 U158 ( .A1(n232), .A2(n57), .B1(n230), .B2(n59), .ZN(n144) );
  AOI221_X1 U159 ( .B1(n53), .B2(n235), .C1(n54), .C2(A[13]), .A(n133), .ZN(
        n45) );
  OAI22_X1 U160 ( .A1(n234), .A2(n57), .B1(n232), .B2(n59), .ZN(n133) );
  AOI222_X1 U161 ( .A1(n12), .A2(n17), .B1(n43), .B2(n146), .C1(n10), .C2(n39), 
        .ZN(n145) );
  OAI221_X1 U162 ( .B1(n46), .B2(n222), .C1(n168), .C2(n221), .A(n151), .ZN(
        n146) );
  OAI221_X1 U163 ( .B1(n20), .B2(n40), .C1(n41), .C2(n180), .A(n42), .ZN(B[3])
         );
  AOI222_X1 U164 ( .A1(n12), .A2(n24), .B1(n43), .B2(n44), .C1(n10), .C2(n23), 
        .ZN(n42) );
  OAI221_X1 U165 ( .B1(n46), .B2(n215), .C1(n168), .C2(n224), .A(n50), .ZN(n44) );
  INV_X1 U166 ( .A(A[19]), .ZN(n120) );
  INV_X1 U167 ( .A(A[30]), .ZN(n111) );
  INV_X1 U168 ( .A(A[31]), .ZN(n213) );
  INV_X1 U169 ( .A(A[29]), .ZN(n113) );
  INV_X1 U170 ( .A(A[18]), .ZN(n136) );
  INV_X1 U171 ( .A(A[11]), .ZN(n232) );
  INV_X1 U172 ( .A(A[23]), .ZN(n208) );
  INV_X1 U173 ( .A(A[21]), .ZN(n206) );
  INV_X1 U174 ( .A(A[28]), .ZN(n114) );
  INV_X1 U175 ( .A(A[16]), .ZN(n202) );
  INV_X1 U176 ( .A(A[17]), .ZN(n203) );
  INV_X1 U177 ( .A(A[27]), .ZN(n212) );
  INV_X1 U178 ( .A(A[10]), .ZN(n230) );
  INV_X1 U179 ( .A(A[9]), .ZN(n228) );
  AOI221_X1 U180 ( .B1(n53), .B2(n225), .C1(n54), .C2(A[7]), .A(n90), .ZN(n32)
         );
  OAI22_X1 U181 ( .A1(n215), .A2(n57), .B1(n224), .B2(n59), .ZN(n90) );
  CLKBUF_X1 U182 ( .A(SH[4]), .Z(n178) );
  AOI22_X1 U183 ( .A1(A[1]), .A2(n166), .B1(A[0]), .B2(n164), .ZN(n151) );
  AOI22_X1 U184 ( .A1(n220), .A2(n166), .B1(A[1]), .B2(n164), .ZN(n89) );
  INV_X1 U185 ( .A(A[8]), .ZN(n226) );
  AOI22_X1 U186 ( .A1(A[3]), .A2(n166), .B1(n220), .B2(n164), .ZN(n67) );
  AOI22_X1 U187 ( .A1(A[4]), .A2(n166), .B1(A[3]), .B2(n164), .ZN(n50) );
  NAND2_X1 U188 ( .A1(SH[1]), .A2(n217), .ZN(n48) );
  NOR2_X1 U189 ( .A1(SH[0]), .A2(SH[1]), .ZN(n52) );
  NOR2_X1 U190 ( .A1(n217), .A2(SH[1]), .ZN(n51) );
  NAND2_X1 U191 ( .A1(SH[1]), .A2(SH[0]), .ZN(n46) );
  NOR2_X1 U192 ( .A1(n219), .A2(SH[2]), .ZN(n78) );
  AND2_X1 U193 ( .A1(SH[2]), .A2(n148), .ZN(n12) );
  INV_X1 U194 ( .A(A[7]), .ZN(n214) );
  INV_X1 U195 ( .A(A[6]), .ZN(n215) );
  INV_X1 U196 ( .A(A[15]), .ZN(n216) );
  INV_X1 U197 ( .A(SH[0]), .ZN(n217) );
  INV_X1 U198 ( .A(SH[2]), .ZN(n218) );
  INV_X1 U199 ( .A(n221), .ZN(n220) );
  INV_X1 U200 ( .A(A[2]), .ZN(n221) );
  INV_X1 U201 ( .A(A[3]), .ZN(n222) );
  INV_X1 U202 ( .A(A[4]), .ZN(n223) );
  INV_X1 U203 ( .A(A[5]), .ZN(n224) );
  INV_X1 U204 ( .A(n226), .ZN(n225) );
  INV_X1 U205 ( .A(n228), .ZN(n227) );
  INV_X1 U206 ( .A(n230), .ZN(n229) );
  INV_X1 U207 ( .A(n232), .ZN(n231) );
  INV_X1 U208 ( .A(n234), .ZN(n233) );
  INV_X1 U209 ( .A(A[12]), .ZN(n234) );
  INV_X1 U210 ( .A(n236), .ZN(n235) );
  INV_X1 U211 ( .A(A[14]), .ZN(n236) );
  INV_X1 U212 ( .A(A[20]), .ZN(n237) );
  INV_X1 U213 ( .A(A[24]), .ZN(n238) );
  INV_X1 U214 ( .A(A[25]), .ZN(n239) );
  INV_X1 U215 ( .A(A[26]), .ZN(n240) );
endmodule


module SHIFTER_GENERIC_N32_DW_sla_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n117, n118, n119, n121, n122, n123, n126, n128,
         n129, n130, n131, n132, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n145, n147, n150, n151, n152, n155, n157, n159, n160,
         n161, n162, n164, n166, n167, n168, n170, n171, n172, n174, n180,
         n181, n185, n186, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230;

  MUX2_X1 U142 ( .A(A[1]), .B(B[0]), .S(n35), .Z(n80) );
  CLKBUF_X3 U2 ( .A(n180), .Z(n185) );
  BUF_X2 U3 ( .A(n180), .Z(n186) );
  INV_X2 U4 ( .A(n186), .ZN(n181) );
  NOR2_X1 U5 ( .A1(n215), .A2(SH[3]), .ZN(n74) );
  INV_X1 U6 ( .A(n12), .ZN(n59) );
  INV_X1 U7 ( .A(n4), .ZN(n130) );
  NAND2_X1 U8 ( .A1(n186), .A2(B[0]), .ZN(n4) );
  INV_X1 U9 ( .A(n35), .ZN(n27) );
  AOI221_X1 U10 ( .B1(n102), .B2(n74), .C1(n103), .C2(n174), .A(n89), .ZN(n7)
         );
  AOI221_X1 U11 ( .B1(n80), .B2(n74), .C1(n73), .C2(n174), .A(n89), .ZN(n8) );
  NAND2_X1 U12 ( .A1(n74), .A2(n181), .ZN(n12) );
  AOI21_X1 U13 ( .B1(n102), .B2(n174), .A(n114), .ZN(n40) );
  AOI21_X1 U14 ( .B1(n95), .B2(n174), .A(n114), .ZN(n10) );
  AOI21_X1 U15 ( .B1(n87), .B2(n174), .A(n114), .ZN(n9) );
  INV_X1 U16 ( .A(n56), .ZN(n17) );
  OAI21_X1 U17 ( .B1(n185), .B2(n29), .A(n4), .ZN(B[14]) );
  OAI21_X1 U18 ( .B1(n185), .B2(n13), .A(n4), .ZN(B[15]) );
  OAI21_X1 U19 ( .B1(n185), .B2(n42), .A(n4), .ZN(B[13]) );
  OAI21_X1 U20 ( .B1(n185), .B2(n64), .A(n4), .ZN(B[10]) );
  OAI21_X1 U21 ( .B1(n185), .B2(n57), .A(n4), .ZN(B[11]) );
  OAI21_X1 U22 ( .B1(n185), .B2(n49), .A(n4), .ZN(B[12]) );
  OAI21_X1 U23 ( .B1(n185), .B2(n6), .A(n4), .ZN(B[7]) );
  OAI21_X1 U24 ( .B1(n185), .B2(n5), .A(n4), .ZN(B[8]) );
  OAI21_X1 U25 ( .B1(n185), .B2(n3), .A(n4), .ZN(B[9]) );
  INV_X1 U26 ( .A(n108), .ZN(n89) );
  INV_X1 U27 ( .A(n107), .ZN(n44) );
  OAI21_X1 U28 ( .B1(n185), .B2(n40), .A(n4), .ZN(B[2]) );
  OAI21_X1 U29 ( .B1(n185), .B2(n117), .A(n4), .ZN(B[1]) );
  OAI21_X1 U30 ( .B1(n185), .B2(n9), .A(n4), .ZN(B[4]) );
  OAI21_X1 U31 ( .B1(n185), .B2(n8), .A(n4), .ZN(B[5]) );
  OAI21_X1 U32 ( .B1(n185), .B2(n7), .A(n4), .ZN(B[6]) );
  AOI21_X1 U33 ( .B1(n80), .B2(n174), .A(n114), .ZN(n117) );
  INV_X1 U34 ( .A(n21), .ZN(n38) );
  INV_X1 U35 ( .A(n23), .ZN(n39) );
  OAI222_X1 U36 ( .A1(n35), .A2(n220), .B1(n218), .B2(n34), .C1(n217), .C2(
        n214), .ZN(n102) );
  INV_X1 U37 ( .A(n34), .ZN(n26) );
  OAI221_X1 U38 ( .B1(n34), .B2(n222), .C1(n35), .C2(n223), .A(n145), .ZN(n73)
         );
  OAI221_X1 U39 ( .B1(n218), .B2(n21), .C1(n217), .C2(n23), .A(n162), .ZN(n95)
         );
  OAI221_X1 U40 ( .B1(n21), .B2(n220), .C1(n218), .C2(n23), .A(n155), .ZN(n87)
         );
  NAND2_X1 U41 ( .A1(n76), .A2(n181), .ZN(n56) );
  AOI221_X1 U42 ( .B1(n26), .B2(n204), .C1(n27), .C2(n206), .A(n126), .ZN(n107) );
  OAI22_X1 U43 ( .A1(n212), .A2(n21), .B1(n230), .B2(n23), .ZN(n126) );
  AOI221_X1 U44 ( .B1(n95), .B2(n74), .C1(n96), .C2(n174), .A(n89), .ZN(n6) );
  AOI221_X1 U45 ( .B1(n87), .B2(n74), .C1(n88), .C2(n174), .A(n89), .ZN(n5) );
  AOI221_X1 U46 ( .B1(n96), .B2(n74), .C1(n93), .C2(n174), .A(n160), .ZN(n57)
         );
  INV_X1 U47 ( .A(n161), .ZN(n160) );
  AOI21_X1 U48 ( .B1(n79), .B2(n95), .A(n81), .ZN(n161) );
  AOI221_X1 U49 ( .B1(n88), .B2(n74), .C1(n85), .C2(n174), .A(n151), .ZN(n49)
         );
  INV_X1 U50 ( .A(n152), .ZN(n151) );
  AOI21_X1 U51 ( .B1(n79), .B2(n87), .A(n81), .ZN(n152) );
  AOI221_X1 U52 ( .B1(n100), .B2(n74), .C1(n66), .C2(n174), .A(n138), .ZN(n29)
         );
  INV_X1 U53 ( .A(n139), .ZN(n138) );
  AOI22_X1 U54 ( .A1(n136), .A2(n102), .B1(n79), .B2(n103), .ZN(n139) );
  AOI221_X1 U55 ( .B1(n75), .B2(n74), .C1(n71), .C2(n174), .A(n141), .ZN(n42)
         );
  INV_X1 U56 ( .A(n142), .ZN(n141) );
  AOI22_X1 U57 ( .A1(n136), .A2(n80), .B1(n79), .B2(n73), .ZN(n142) );
  AOI221_X1 U58 ( .B1(n73), .B2(n74), .C1(n75), .C2(n174), .A(n77), .ZN(n3) );
  INV_X1 U59 ( .A(n78), .ZN(n77) );
  AOI21_X1 U60 ( .B1(n79), .B2(n80), .A(n81), .ZN(n78) );
  AOI221_X1 U61 ( .B1(n103), .B2(n74), .C1(n100), .C2(n174), .A(n167), .ZN(n64) );
  INV_X1 U62 ( .A(n168), .ZN(n167) );
  AOI21_X1 U63 ( .B1(n79), .B2(n102), .A(n81), .ZN(n168) );
  AOI222_X1 U64 ( .A1(n59), .A2(n31), .B1(n19), .B2(n66), .C1(n15), .C2(n100), 
        .ZN(n99) );
  AOI222_X1 U65 ( .A1(n59), .A2(n44), .B1(n19), .B2(n71), .C1(n15), .C2(n75), 
        .ZN(n106) );
  AOI222_X1 U66 ( .A1(n59), .A2(n51), .B1(n19), .B2(n85), .C1(n15), .C2(n88), 
        .ZN(n112) );
  AOI222_X1 U67 ( .A1(n59), .A2(n16), .B1(n19), .B2(n60), .C1(n15), .C2(n93), 
        .ZN(n92) );
  AOI222_X1 U68 ( .A1(n59), .A2(n60), .B1(n19), .B2(n93), .C1(n15), .C2(n96), 
        .ZN(n118) );
  AOI222_X1 U69 ( .A1(n59), .A2(n46), .B1(n19), .B2(n44), .C1(n15), .C2(n71), 
        .ZN(n70) );
  AOI222_X1 U70 ( .A1(n59), .A2(n53), .B1(n19), .B2(n51), .C1(n15), .C2(n85), 
        .ZN(n84) );
  OAI221_X1 U71 ( .B1(n72), .B2(n56), .C1(n8), .C2(n181), .A(n106), .ZN(B[21])
         );
  OAI221_X1 U72 ( .B1(n67), .B2(n56), .C1(n7), .C2(n181), .A(n99), .ZN(B[22])
         );
  OAI221_X1 U73 ( .B1(n94), .B2(n56), .C1(n10), .C2(n181), .A(n118), .ZN(B[19]) );
  OAI21_X1 U74 ( .B1(n217), .B2(n215), .A(n108), .ZN(n114) );
  NOR2_X1 U75 ( .A1(n215), .A2(n108), .ZN(n81) );
  NAND2_X1 U76 ( .A1(n213), .A2(n214), .ZN(n35) );
  BUF_X1 U77 ( .A(n76), .Z(n174) );
  AND2_X1 U78 ( .A1(n131), .A2(n215), .ZN(n19) );
  OAI221_X1 U79 ( .B1(n107), .B2(n56), .C1(n117), .C2(n181), .A(n123), .ZN(
        B[17]) );
  AOI222_X1 U80 ( .A1(n59), .A2(n71), .B1(n19), .B2(n75), .C1(n15), .C2(n73), 
        .ZN(n123) );
  AND2_X1 U81 ( .A1(SH[3]), .A2(n215), .ZN(n79) );
  NAND2_X1 U82 ( .A1(SH[3]), .A2(B[0]), .ZN(n108) );
  INV_X1 U83 ( .A(n171), .ZN(n103) );
  AOI221_X1 U84 ( .B1(n38), .B2(n221), .C1(A[3]), .C2(n39), .A(n172), .ZN(n171) );
  OAI22_X1 U85 ( .A1(n223), .A2(n34), .B1(n211), .B2(n35), .ZN(n172) );
  INV_X1 U86 ( .A(n94), .ZN(n16) );
  INV_X1 U87 ( .A(n101), .ZN(n31) );
  INV_X1 U88 ( .A(n113), .ZN(n51) );
  OAI221_X1 U89 ( .B1(n86), .B2(n56), .C1(n9), .C2(n181), .A(n112), .ZN(B[20])
         );
  INV_X1 U90 ( .A(n61), .ZN(n20) );
  INV_X1 U91 ( .A(n72), .ZN(n46) );
  INV_X1 U92 ( .A(n67), .ZN(n33) );
  INV_X1 U93 ( .A(n86), .ZN(n53) );
  INV_X1 U94 ( .A(n205), .ZN(n204) );
  INV_X1 U95 ( .A(n207), .ZN(n206) );
  OAI221_X1 U96 ( .B1(n11), .B2(n56), .C1(n57), .C2(n181), .A(n58), .ZN(B[27])
         );
  AOI222_X1 U97 ( .A1(n59), .A2(n20), .B1(n19), .B2(n16), .C1(n15), .C2(n60), 
        .ZN(n58) );
  OAI221_X1 U98 ( .B1(n28), .B2(n56), .C1(n64), .C2(n181), .A(n65), .ZN(B[26])
         );
  AOI222_X1 U99 ( .A1(n59), .A2(n33), .B1(n19), .B2(n31), .C1(n15), .C2(n66), 
        .ZN(n65) );
  OAI221_X1 U100 ( .B1(n11), .B2(n12), .C1(n13), .C2(n181), .A(n14), .ZN(B[31]) );
  AOI222_X1 U101 ( .A1(n15), .A2(n16), .B1(n17), .B2(n18), .C1(n19), .C2(n20), 
        .ZN(n14) );
  OAI221_X1 U102 ( .B1(n21), .B2(n22), .C1(n23), .C2(n24), .A(n25), .ZN(n18)
         );
  OAI221_X1 U103 ( .B1(n48), .B2(n12), .C1(n49), .C2(n181), .A(n50), .ZN(B[28]) );
  AOI222_X1 U104 ( .A1(n15), .A2(n51), .B1(n17), .B2(n52), .C1(n19), .C2(n53), 
        .ZN(n50) );
  OAI221_X1 U105 ( .B1(n34), .B2(n209), .C1(n35), .C2(n24), .A(n55), .ZN(n52)
         );
  OAI221_X1 U106 ( .B1(n28), .B2(n12), .C1(n29), .C2(n181), .A(n30), .ZN(B[30]) );
  AOI222_X1 U107 ( .A1(n15), .A2(n31), .B1(n17), .B2(n32), .C1(n19), .C2(n33), 
        .ZN(n30) );
  OAI221_X1 U108 ( .B1(n34), .B2(n22), .C1(n35), .C2(n36), .A(n37), .ZN(n32)
         );
  OAI221_X1 U109 ( .B1(n41), .B2(n12), .C1(n42), .C2(n181), .A(n43), .ZN(B[29]) );
  AOI222_X1 U110 ( .A1(n15), .A2(n44), .B1(n17), .B2(n45), .C1(n19), .C2(n46), 
        .ZN(n43) );
  OAI221_X1 U111 ( .B1(n34), .B2(n24), .C1(n35), .C2(n22), .A(n47), .ZN(n45)
         );
  OAI221_X1 U112 ( .B1(n101), .B2(n56), .C1(n40), .C2(n181), .A(n121), .ZN(
        B[18]) );
  AOI222_X1 U113 ( .A1(n59), .A2(n66), .B1(n19), .B2(n100), .C1(n15), .C2(n103), .ZN(n121) );
  OAI221_X1 U114 ( .B1(n128), .B2(n12), .C1(n113), .C2(n56), .A(n129), .ZN(
        B[16]) );
  INV_X1 U115 ( .A(n85), .ZN(n128) );
  AOI221_X1 U116 ( .B1(n15), .B2(n87), .C1(n19), .C2(n88), .A(n130), .ZN(n129)
         );
  AND2_X1 U117 ( .A1(SH[3]), .A2(n181), .ZN(n131) );
  OAI21_X1 U118 ( .B1(n185), .B2(n10), .A(n4), .ZN(B[3]) );
  AOI221_X1 U119 ( .B1(n93), .B2(n74), .C1(n60), .C2(n174), .A(n134), .ZN(n13)
         );
  INV_X1 U120 ( .A(n135), .ZN(n134) );
  AOI22_X1 U121 ( .A1(n136), .A2(n95), .B1(n79), .B2(n96), .ZN(n135) );
  OAI221_X1 U122 ( .B1(n61), .B2(n56), .C1(n6), .C2(n181), .A(n92), .ZN(B[23])
         );
  INV_X1 U123 ( .A(n209), .ZN(n208) );
  OAI221_X1 U124 ( .B1(n34), .B2(n210), .C1(n35), .C2(n224), .A(n159), .ZN(n88) );
  OAI221_X1 U125 ( .B1(n34), .B2(n211), .C1(n35), .C2(n210), .A(n166), .ZN(n96) );
  OAI221_X1 U126 ( .B1(n34), .B2(n227), .C1(n35), .C2(n228), .A(n157), .ZN(n85) );
  AOI22_X1 U127 ( .A1(A[10]), .A2(n38), .B1(A[9]), .B2(n39), .ZN(n157) );
  OAI221_X1 U128 ( .B1(n34), .B2(n226), .C1(n35), .C2(n227), .A(n164), .ZN(n93) );
  OAI221_X1 U129 ( .B1(n34), .B2(n224), .C1(n35), .C2(n225), .A(n150), .ZN(n75) );
  OAI221_X1 U130 ( .B1(n34), .B2(n225), .C1(n35), .C2(n226), .A(n170), .ZN(
        n100) );
  OAI221_X1 U131 ( .B1(n34), .B2(n228), .C1(n35), .C2(n229), .A(n147), .ZN(n71) );
  AOI22_X1 U132 ( .A1(A[11]), .A2(n38), .B1(A[10]), .B2(n39), .ZN(n147) );
  OAI221_X1 U133 ( .B1(n34), .B2(n229), .C1(n35), .C2(n230), .A(n140), .ZN(n66) );
  AOI22_X1 U134 ( .A1(A[12]), .A2(n38), .B1(A[11]), .B2(n39), .ZN(n140) );
  OAI221_X1 U135 ( .B1(n34), .B2(n230), .C1(n35), .C2(n212), .A(n137), .ZN(n60) );
  AOI22_X1 U136 ( .A1(A[13]), .A2(n38), .B1(A[12]), .B2(n39), .ZN(n137) );
  AOI221_X1 U137 ( .B1(n26), .B2(A[24]), .C1(n27), .C2(A[25]), .A(n82), .ZN(
        n41) );
  INV_X1 U138 ( .A(n83), .ZN(n82) );
  AOI22_X1 U139 ( .A1(A[23]), .A2(n38), .B1(A[22]), .B2(n39), .ZN(n83) );
  AOI221_X1 U140 ( .B1(n26), .B2(A[23]), .C1(n27), .C2(A[24]), .A(n90), .ZN(
        n48) );
  INV_X1 U141 ( .A(n91), .ZN(n90) );
  AOI22_X1 U143 ( .A1(A[22]), .A2(n38), .B1(A[21]), .B2(n39), .ZN(n91) );
  AOI221_X1 U144 ( .B1(n26), .B2(A[25]), .C1(n27), .C2(A[26]), .A(n68), .ZN(
        n28) );
  INV_X1 U145 ( .A(n69), .ZN(n68) );
  AOI22_X1 U146 ( .A1(A[24]), .A2(n38), .B1(A[23]), .B2(n39), .ZN(n69) );
  AOI221_X1 U147 ( .B1(n26), .B2(A[26]), .C1(n27), .C2(n208), .A(n62), .ZN(n11) );
  INV_X1 U148 ( .A(n63), .ZN(n62) );
  AOI22_X1 U149 ( .A1(A[25]), .A2(n38), .B1(A[24]), .B2(n39), .ZN(n63) );
  AOI221_X1 U150 ( .B1(n26), .B2(A[22]), .C1(n27), .C2(A[23]), .A(n97), .ZN(
        n61) );
  INV_X1 U151 ( .A(n98), .ZN(n97) );
  AOI22_X1 U152 ( .A1(A[21]), .A2(n38), .B1(A[20]), .B2(n39), .ZN(n98) );
  AOI221_X1 U153 ( .B1(n26), .B2(A[20]), .C1(n27), .C2(A[21]), .A(n109), .ZN(
        n72) );
  OAI22_X1 U154 ( .A1(n110), .A2(n21), .B1(n111), .B2(n23), .ZN(n109) );
  INV_X1 U155 ( .A(A[19]), .ZN(n110) );
  AOI221_X1 U156 ( .B1(n26), .B2(A[21]), .C1(n27), .C2(A[22]), .A(n104), .ZN(
        n67) );
  INV_X1 U157 ( .A(n105), .ZN(n104) );
  AOI22_X1 U158 ( .A1(A[20]), .A2(n38), .B1(A[19]), .B2(n39), .ZN(n105) );
  AOI221_X1 U159 ( .B1(n26), .B2(A[18]), .C1(n27), .C2(A[19]), .A(n119), .ZN(
        n94) );
  OAI22_X1 U160 ( .A1(n207), .A2(n21), .B1(n205), .B2(n23), .ZN(n119) );
  AOI221_X1 U161 ( .B1(n26), .B2(n206), .C1(n27), .C2(A[18]), .A(n122), .ZN(
        n101) );
  OAI22_X1 U162 ( .A1(n205), .A2(n21), .B1(n212), .B2(n23), .ZN(n122) );
  AOI221_X1 U163 ( .B1(n26), .B2(A[19]), .C1(n27), .C2(A[20]), .A(n115), .ZN(
        n86) );
  OAI22_X1 U164 ( .A1(n111), .A2(n21), .B1(n207), .B2(n23), .ZN(n115) );
  AOI221_X1 U165 ( .B1(n26), .B2(A[15]), .C1(n27), .C2(n204), .A(n132), .ZN(
        n113) );
  OAI22_X1 U166 ( .A1(n230), .A2(n21), .B1(n229), .B2(n23), .ZN(n132) );
  OAI221_X1 U167 ( .B1(n48), .B2(n56), .C1(n5), .C2(n181), .A(n84), .ZN(B[24])
         );
  OAI221_X1 U168 ( .B1(n41), .B2(n56), .C1(n3), .C2(n181), .A(n70), .ZN(B[25])
         );
  AOI22_X1 U169 ( .A1(A[30]), .A2(n26), .B1(A[31]), .B2(n27), .ZN(n25) );
  AOI22_X1 U170 ( .A1(A[28]), .A2(n38), .B1(n208), .B2(n39), .ZN(n37) );
  AOI22_X1 U171 ( .A1(A[26]), .A2(n38), .B1(A[25]), .B2(n39), .ZN(n55) );
  AOI22_X1 U172 ( .A1(n208), .A2(n38), .B1(A[26]), .B2(n39), .ZN(n47) );
  INV_X1 U173 ( .A(A[16]), .ZN(n205) );
  INV_X1 U174 ( .A(A[17]), .ZN(n207) );
  INV_X1 U175 ( .A(A[18]), .ZN(n111) );
  CLKBUF_X1 U176 ( .A(SH[4]), .Z(n180) );
  INV_X1 U177 ( .A(A[28]), .ZN(n24) );
  INV_X1 U178 ( .A(A[29]), .ZN(n22) );
  INV_X1 U179 ( .A(A[27]), .ZN(n209) );
  INV_X1 U180 ( .A(A[30]), .ZN(n36) );
  INV_X1 U181 ( .A(A[2]), .ZN(n220) );
  AOI22_X1 U182 ( .A1(A[9]), .A2(n38), .B1(A[8]), .B2(n39), .ZN(n164) );
  AOI22_X1 U183 ( .A1(A[3]), .A2(n38), .B1(n219), .B2(n39), .ZN(n145) );
  AOI22_X1 U184 ( .A1(n26), .A2(A[3]), .B1(n221), .B2(n27), .ZN(n155) );
  AOI22_X1 U185 ( .A1(n26), .A2(n219), .B1(A[3]), .B2(n27), .ZN(n162) );
  AOI22_X1 U186 ( .A1(A[6]), .A2(n38), .B1(A[5]), .B2(n39), .ZN(n159) );
  AOI22_X1 U187 ( .A1(A[5]), .A2(n38), .B1(n221), .B2(n39), .ZN(n166) );
  NAND2_X1 U188 ( .A1(SH[0]), .A2(n214), .ZN(n34) );
  AOI22_X1 U189 ( .A1(A[7]), .A2(n38), .B1(A[6]), .B2(n39), .ZN(n150) );
  AOI22_X1 U190 ( .A1(A[8]), .A2(n38), .B1(A[7]), .B2(n39), .ZN(n170) );
  NAND2_X1 U191 ( .A1(SH[1]), .A2(n213), .ZN(n21) );
  NAND2_X1 U192 ( .A1(SH[0]), .A2(SH[1]), .ZN(n23) );
  AND2_X1 U193 ( .A1(SH[2]), .A2(SH[3]), .ZN(n136) );
  AND2_X1 U194 ( .A1(n131), .A2(SH[2]), .ZN(n15) );
  NOR2_X1 U195 ( .A1(SH[2]), .A2(SH[3]), .ZN(n76) );
  INV_X1 U196 ( .A(A[7]), .ZN(n210) );
  INV_X1 U197 ( .A(A[6]), .ZN(n211) );
  INV_X1 U198 ( .A(A[15]), .ZN(n212) );
  INV_X1 U199 ( .A(SH[0]), .ZN(n213) );
  INV_X1 U200 ( .A(SH[1]), .ZN(n214) );
  INV_X1 U201 ( .A(SH[2]), .ZN(n215) );
  INV_X1 U202 ( .A(n217), .ZN(B[0]) );
  INV_X1 U203 ( .A(A[0]), .ZN(n217) );
  INV_X1 U204 ( .A(A[1]), .ZN(n218) );
  INV_X1 U205 ( .A(n220), .ZN(n219) );
  INV_X1 U206 ( .A(n222), .ZN(n221) );
  INV_X1 U207 ( .A(A[4]), .ZN(n222) );
  INV_X1 U208 ( .A(A[5]), .ZN(n223) );
  INV_X1 U209 ( .A(A[8]), .ZN(n224) );
  INV_X1 U210 ( .A(A[9]), .ZN(n225) );
  INV_X1 U211 ( .A(A[10]), .ZN(n226) );
  INV_X1 U212 ( .A(A[11]), .ZN(n227) );
  INV_X1 U213 ( .A(A[12]), .ZN(n228) );
  INV_X1 U214 ( .A(A[13]), .ZN(n229) );
  INV_X1 U215 ( .A(A[14]), .ZN(n230) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n3,
         n4, n5, n6, n7, n8, n9, n10, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n27), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n27), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n27), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n27), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n27), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n28), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n28), .Z(B[25]) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n28), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n28), .Z(B[23]) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n28), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n28), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n28), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n28), .Z(B[19]) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n28), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n28), .Z(B[17]) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n27), .Z(B[16]) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n39), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n39), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n39), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n39), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n39), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n39), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n39), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n39), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n39), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n39), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n39), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n39), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n38), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n38), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n38), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n38), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n38), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n38), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n38), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n38), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n38), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n38), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n38), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n38), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n35), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n35), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n35), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n35), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n35), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n35), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n35), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n35), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n35), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n35), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n35), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n35), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n35), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n35), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n35), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n35), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n36), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n36), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n36), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n36), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n36), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n36), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n36), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n36), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n36), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n36), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n36), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n36), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n33), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n33), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n33), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n33), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n33), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n33), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n32), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n32), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n32), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n32), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n32), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n32), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n32), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n32), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n32), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n32), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n32), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n32), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n31), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n31), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n31), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n31), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n31), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n31), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n31), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n31), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n31), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n31), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n31), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n31), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  INV_X2 U3 ( .A(n37), .ZN(n35) );
  AND2_X1 U4 ( .A1(\ML_int[4][8] ), .A2(n29), .ZN(B[8]) );
  AND2_X1 U5 ( .A1(\ML_int[4][9] ), .A2(n29), .ZN(B[9]) );
  AND2_X1 U6 ( .A1(\ML_int[4][10] ), .A2(n29), .ZN(B[10]) );
  AND2_X1 U7 ( .A1(\ML_int[4][11] ), .A2(n29), .ZN(B[11]) );
  AND2_X1 U8 ( .A1(\ML_int[4][12] ), .A2(n29), .ZN(B[12]) );
  AND2_X1 U9 ( .A1(\ML_int[4][13] ), .A2(n29), .ZN(B[13]) );
  AND2_X1 U10 ( .A1(\ML_int[4][14] ), .A2(n29), .ZN(B[14]) );
  AND2_X1 U11 ( .A1(\ML_int[4][15] ), .A2(n29), .ZN(B[15]) );
  NAND2_X1 U12 ( .A1(\ML_int[3][7] ), .A2(n40), .ZN(n3) );
  NAND2_X1 U13 ( .A1(\ML_int[3][6] ), .A2(n40), .ZN(n4) );
  NAND2_X1 U14 ( .A1(\ML_int[3][4] ), .A2(n40), .ZN(n6) );
  NAND2_X1 U15 ( .A1(\ML_int[3][5] ), .A2(n40), .ZN(n5) );
  NAND2_X1 U16 ( .A1(\ML_int[3][3] ), .A2(n40), .ZN(n7) );
  NAND2_X1 U17 ( .A1(\ML_int[3][2] ), .A2(n40), .ZN(n8) );
  INV_X1 U18 ( .A(n10), .ZN(\ML_int[4][0] ) );
  INV_X1 U19 ( .A(n6), .ZN(\ML_int[4][4] ) );
  INV_X1 U20 ( .A(n7), .ZN(\ML_int[4][3] ) );
  INV_X1 U21 ( .A(n4), .ZN(\ML_int[4][6] ) );
  INV_X1 U22 ( .A(n5), .ZN(\ML_int[4][5] ) );
  INV_X1 U23 ( .A(n8), .ZN(\ML_int[4][2] ) );
  INV_X1 U24 ( .A(n9), .ZN(\ML_int[4][1] ) );
  INV_X1 U25 ( .A(n3), .ZN(\ML_int[4][7] ) );
  NOR2_X1 U26 ( .A1(n27), .A2(n6), .ZN(B[4]) );
  NOR2_X1 U27 ( .A1(n27), .A2(n5), .ZN(B[5]) );
  NOR2_X1 U28 ( .A1(n27), .A2(n4), .ZN(B[6]) );
  NOR2_X1 U29 ( .A1(n27), .A2(n3), .ZN(B[7]) );
  INV_X1 U30 ( .A(n41), .ZN(n38) );
  INV_X1 U31 ( .A(n41), .ZN(n39) );
  NAND2_X1 U32 ( .A1(\ML_int[3][1] ), .A2(n40), .ZN(n9) );
  NAND2_X1 U33 ( .A1(\ML_int[3][0] ), .A2(n40), .ZN(n10) );
  INV_X1 U34 ( .A(n34), .ZN(n31) );
  AND2_X1 U35 ( .A1(\ML_int[2][3] ), .A2(n37), .ZN(\ML_int[3][3] ) );
  AND2_X1 U36 ( .A1(\ML_int[2][2] ), .A2(n37), .ZN(\ML_int[3][2] ) );
  AND2_X1 U37 ( .A1(\ML_int[2][1] ), .A2(n37), .ZN(\ML_int[3][1] ) );
  AND2_X1 U38 ( .A1(\ML_int[1][1] ), .A2(n34), .ZN(\ML_int[2][1] ) );
  INV_X1 U39 ( .A(n29), .ZN(n27) );
  INV_X1 U40 ( .A(n37), .ZN(n36) );
  INV_X1 U41 ( .A(n34), .ZN(n32) );
  INV_X1 U42 ( .A(n29), .ZN(n28) );
  AND2_X1 U43 ( .A1(\ML_int[2][0] ), .A2(n37), .ZN(\ML_int[3][0] ) );
  AND2_X1 U44 ( .A1(\ML_int[1][0] ), .A2(n34), .ZN(\ML_int[2][0] ) );
  NOR2_X1 U45 ( .A1(n27), .A2(n8), .ZN(B[2]) );
  NOR2_X1 U46 ( .A1(n27), .A2(n7), .ZN(B[3]) );
  NOR2_X1 U47 ( .A1(n27), .A2(n9), .ZN(B[1]) );
  NOR2_X1 U48 ( .A1(n27), .A2(n10), .ZN(B[0]) );
  INV_X1 U49 ( .A(SH[4]), .ZN(n29) );
  AND2_X1 U50 ( .A1(A[0]), .A2(n30), .ZN(\ML_int[1][0] ) );
  INV_X1 U51 ( .A(SH[0]), .ZN(n30) );
  INV_X1 U52 ( .A(SH[2]), .ZN(n37) );
  INV_X1 U53 ( .A(SH[1]), .ZN(n34) );
  INV_X1 U54 ( .A(n34), .ZN(n33) );
  INV_X1 U55 ( .A(SH[3]), .ZN(n40) );
  INV_X1 U56 ( .A(SH[3]), .ZN(n41) );
endmodule


module p4adder_N32_0 ( A, B, Cin, S, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout;

  wire   [8:0] C;

  CarryGen_N32_0 Cgen ( .A(A), .B(B), .Cin(Cin), .C(C) );
  SumGen_N32_0 Sgen ( .A(A), .B(B), .C(C), .S(S), .Cout(Cout) );
endmodule


module xor_gen_N32_1 ( A, B, C );
  input [31:0] A;
  input [31:0] B;
  output [31:0] C;


  XOR2_X1 U1 ( .A(A[2]), .B(B[2]), .Z(C[2]) );
  XOR2_X1 U2 ( .A(A[0]), .B(B[0]), .Z(C[0]) );
  XOR2_X1 U3 ( .A(A[1]), .B(B[1]), .Z(C[1]) );
  XOR2_X1 U4 ( .A(A[31]), .B(B[31]), .Z(C[31]) );
  XOR2_X1 U5 ( .A(A[11]), .B(B[11]), .Z(C[11]) );
  XOR2_X1 U6 ( .A(A[9]), .B(B[9]), .Z(C[9]) );
  XOR2_X1 U7 ( .A(A[13]), .B(B[13]), .Z(C[13]) );
  XOR2_X1 U8 ( .A(A[6]), .B(B[6]), .Z(C[6]) );
  XOR2_X1 U9 ( .A(A[10]), .B(B[10]), .Z(C[10]) );
  XOR2_X1 U10 ( .A(A[14]), .B(B[14]), .Z(C[14]) );
  XOR2_X1 U11 ( .A(A[12]), .B(B[12]), .Z(C[12]) );
  XOR2_X1 U12 ( .A(A[15]), .B(B[15]), .Z(C[15]) );
  XOR2_X1 U13 ( .A(A[17]), .B(B[17]), .Z(C[17]) );
  XOR2_X1 U14 ( .A(A[21]), .B(B[21]), .Z(C[21]) );
  XOR2_X1 U15 ( .A(A[19]), .B(B[19]), .Z(C[19]) );
  XOR2_X1 U16 ( .A(A[23]), .B(B[23]), .Z(C[23]) );
  XOR2_X1 U17 ( .A(A[18]), .B(B[18]), .Z(C[18]) );
  XOR2_X1 U18 ( .A(A[16]), .B(B[16]), .Z(C[16]) );
  XOR2_X1 U19 ( .A(A[25]), .B(B[25]), .Z(C[25]) );
  XOR2_X1 U20 ( .A(A[22]), .B(B[22]), .Z(C[22]) );
  XOR2_X1 U21 ( .A(A[20]), .B(B[20]), .Z(C[20]) );
  XOR2_X1 U22 ( .A(A[27]), .B(B[27]), .Z(C[27]) );
  XOR2_X1 U23 ( .A(A[29]), .B(B[29]), .Z(C[29]) );
  XOR2_X1 U24 ( .A(A[26]), .B(B[26]), .Z(C[26]) );
  XOR2_X1 U25 ( .A(A[28]), .B(B[28]), .Z(C[28]) );
  XOR2_X1 U26 ( .A(A[24]), .B(B[24]), .Z(C[24]) );
  XOR2_X1 U27 ( .A(A[30]), .B(B[30]), .Z(C[30]) );
  XOR2_X1 U28 ( .A(A[3]), .B(B[3]), .Z(C[3]) );
  XOR2_X1 U29 ( .A(A[4]), .B(B[4]), .Z(C[4]) );
  XOR2_X1 U30 ( .A(A[5]), .B(B[5]), .Z(C[5]) );
  XOR2_X1 U31 ( .A(A[7]), .B(B[7]), .Z(C[7]) );
  XOR2_X1 U32 ( .A(A[8]), .B(B[8]), .Z(C[8]) );
endmodule


module MUX21_647 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_647 UIV ( .A(S), .Y(SB) );
  ND2_1941 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_1940 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_1939 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_742 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_742 UIV ( .A(S), .Y(SB) );
  ND2_2226 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2225 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2224 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_743 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_743 UIV ( .A(S), .Y(SB) );
  ND2_2229 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2228 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2227 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_887 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_887 UIV ( .A(S), .Y(SB) );
  ND2_2661 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2660 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2659 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_913 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_913 UIV ( .A(S), .Y(SB) );
  ND2_2739 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2738 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2737 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module IV_942 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module ND2_2827 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module ND2_2828 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(Y) );
endmodule


module ND2_0 ( A, B, Y );
  input A, B;
  output Y;


  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(Y) );
endmodule


module IV_0 ( A, Y );
  input A;
  output Y;


  INV_X1 U1 ( .A(A), .ZN(Y) );
endmodule


module MUX21_GENERIC_N32_9 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_544 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_543 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_542 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_541 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_540 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_539 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_538 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_537 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_536 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_535 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_534 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_533 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_532 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_531 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_530 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_529 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_528 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_527 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_526 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_525 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_524 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_523 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_522 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_521 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_520 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_519 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_518 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_517 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_516 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_515 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_514 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_513 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n5) );
  BUF_X1 U2 ( .A(n3), .Z(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_10 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_576 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_575 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_574 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_573 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_572 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_571 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_570 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_569 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_568 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_567 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_566 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_565 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_564 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_563 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_562 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_561 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_560 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_559 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_558 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_557 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_556 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_555 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_554 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_553 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_552 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_551 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_550 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_549 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_548 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_547 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_546 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_545 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n4) );
  BUF_X1 U2 ( .A(n3), .Z(n5) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module mux81_generic_N32 ( A, B, C, D, E, F, G, H, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [31:0] G;
  input [31:0] H;
  input [2:0] S;
  output [31:0] Y;

  wire   [31:0] ABto2;
  wire   [31:0] CDto2;
  wire   [31:0] EFto2;
  wire   [31:0] GHto2;
  wire   [31:0] ABCDto3;
  wire   [31:0] EFGHto3;

  MUX21_GENERIC_N32_7 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_GENERIC_N32_6 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_GENERIC_N32_5 M13 ( .A(E), .B(F), .S(S[0]), .Y(EFto2) );
  MUX21_GENERIC_N32_4 M14 ( .A(G), .B(H), .S(S[0]), .Y(GHto2) );
  MUX21_GENERIC_N32_3 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(ABCDto3) );
  MUX21_GENERIC_N32_2 M22 ( .A(EFto2), .B(GHto2), .S(S[1]), .Y(EFGHto3) );
  MUX21_GENERIC_N32_1 M31 ( .A(ABCDto3), .B(EFGHto3), .S(S[2]), .Y(Y) );
endmodule


module MUX21_GENERIC_N32_11 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_608 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_607 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_606 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_605 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_604 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_603 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_602 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_601 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_600 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_599 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_598 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_597 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_596 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_595 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_594 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_593 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_592 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_591 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_590 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_589 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_588 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_587 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_586 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_585 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_584 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_583 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_582 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_581 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_580 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_579 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_578 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_577 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n4) );
  BUF_X1 U2 ( .A(n3), .Z(n5) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module mux81_logic ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   ABto2, CDto2, EFto2, GHto2, ABCDto3, EFGHto3;

  MUX21_615 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_614 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_613 M13 ( .A(E), .B(F), .S(S[0]), .Y(EFto2) );
  MUX21_612 M14 ( .A(G), .B(H), .S(S[0]), .Y(GHto2) );
  MUX21_611 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(ABCDto3) );
  MUX21_610 M22 ( .A(EFto2), .B(GHto2), .S(S[1]), .Y(EFGHto3) );
  MUX21_609 M31 ( .A(ABCDto3), .B(EFGHto3), .S(S[2]), .Y(Y) );
endmodule


module Boothmul_N16 ( A, B, P );
  input [15:0] A;
  input [15:0] B;
  output [31:0] P;
  wire   \MinusAExt1[5][31] , \MinusAExt1[5][30] , \MinusAExt1[5][29] ,
         \MinusAExt1[5][28] , \MinusAExt1[5][27] , \MinusAExt1[5][26] ,
         \MinusAExt1[5][25] , \MinusAExt1[5][24] , \MinusAExt1[5][23] ,
         \MinusAExt1[5][22] , \MinusAExt1[5][21] , \MinusAExt1[5][20] ,
         \MinusAExt1[5][19] , \MinusAExt1[5][18] , \MinusAExt1[5][17] ,
         \MinusAExt1[5][16] , \MinusAExt1[5][15] , \MinusAExt1[5][14] ,
         \MinusAExt1[5][13] , \MinusAExt1[5][12] , \MinusAExt1[5][11] ,
         \MinusAExt1[5][10] , \MinusAExt2[4][31] , \MinusAExt2[4][30] ,
         \MinusAExt2[4][29] , \MinusAExt2[4][28] , \MinusAExt2[4][27] ,
         \MinusAExt2[4][26] , \MinusAExt2[4][25] , \MinusAExt2[4][24] ,
         \MinusAExt2[4][23] , \MinusAExt2[4][22] , \MinusAExt2[4][21] ,
         \MinusAExt2[4][20] , \MinusAExt2[4][19] , \MinusAExt2[4][18] ,
         \MinusAExt2[4][17] , \MinusAExt2[4][16] , \MinusAExt2[4][15] ,
         \MinusAExt2[4][14] , \MinusAExt2[4][13] , \MinusAExt2[4][12] ,
         \MinusAExt2[4][11] , \MinusAExt2[4][10] , \MinusAExt2[4][9] ,
         \Sel[7][2] , \Sel[7][1] , \Sel[7][0] , \Sel[6][2] , \Sel[6][1] ,
         \Sel[6][0] , \Sel[5][2] , \Sel[5][1] , \Sel[5][0] , \Sel[4][2] ,
         \Sel[4][1] , \Sel[4][0] , \Sel[3][2] , \Sel[3][1] , \Sel[3][0] ,
         \Sel[2][2] , \Sel[2][1] , \Sel[2][0] , \Sel[1][2] , \Sel[1][1] ,
         \Sel[1][0] , \Sel[0][2] , \Sel[0][0] , \Sum[7][31] , \Sum[7][30] ,
         \Sum[7][29] , \Sum[7][28] , \Sum[7][27] , \Sum[7][26] , \Sum[7][25] ,
         \Sum[7][24] , \Sum[7][23] , \Sum[7][22] , \Sum[7][21] , \Sum[7][20] ,
         \Sum[7][19] , \Sum[7][18] , \Sum[7][17] , \Sum[7][16] , \Sum[7][15] ,
         \Sum[7][14] , \Sum[7][13] , \Sum[7][12] , \Sum[7][11] , \Sum[7][10] ,
         \Sum[7][9] , \Sum[7][8] , \Sum[7][7] , \Sum[7][6] , \Sum[7][5] ,
         \Sum[7][4] , \Sum[7][3] , \Sum[7][2] , \Sum[7][1] , \Sum[7][0] ,
         \Sum[6][31] , \Sum[6][30] , \Sum[6][29] , \Sum[6][28] , \Sum[6][27] ,
         \Sum[6][26] , \Sum[6][25] , \Sum[6][24] , \Sum[6][23] , \Sum[6][22] ,
         \Sum[6][21] , \Sum[6][20] , \Sum[6][19] , \Sum[6][18] , \Sum[6][17] ,
         \Sum[6][16] , \Sum[6][15] , \Sum[6][14] , \Sum[6][13] , \Sum[6][12] ,
         \Sum[6][11] , \Sum[6][10] , \Sum[6][9] , \Sum[6][8] , \Sum[6][7] ,
         \Sum[6][6] , \Sum[6][5] , \Sum[6][4] , \Sum[6][3] , \Sum[6][2] ,
         \Sum[6][1] , \Sum[6][0] , \Sum[5][31] , \Sum[5][30] , \Sum[5][29] ,
         \Sum[5][28] , \Sum[5][27] , \Sum[5][26] , \Sum[5][25] , \Sum[5][24] ,
         \Sum[5][23] , \Sum[5][22] , \Sum[5][21] , \Sum[5][20] , \Sum[5][19] ,
         \Sum[5][18] , \Sum[5][17] , \Sum[5][16] , \Sum[5][15] , \Sum[5][14] ,
         \Sum[5][13] , \Sum[5][12] , \Sum[5][11] , \Sum[5][10] , \Sum[5][9] ,
         \Sum[5][8] , \Sum[5][7] , \Sum[5][6] , \Sum[5][5] , \Sum[5][4] ,
         \Sum[5][3] , \Sum[5][2] , \Sum[5][1] , \Sum[5][0] , \Sum[4][31] ,
         \Sum[4][30] , \Sum[4][29] , \Sum[4][28] , \Sum[4][27] , \Sum[4][26] ,
         \Sum[4][25] , \Sum[4][24] , \Sum[4][23] , \Sum[4][22] , \Sum[4][21] ,
         \Sum[4][20] , \Sum[4][19] , \Sum[4][18] , \Sum[4][17] , \Sum[4][16] ,
         \Sum[4][15] , \Sum[4][14] , \Sum[4][13] , \Sum[4][12] , \Sum[4][11] ,
         \Sum[4][10] , \Sum[4][9] , \Sum[4][8] , \Sum[4][7] , \Sum[4][6] ,
         \Sum[4][5] , \Sum[4][4] , \Sum[4][3] , \Sum[4][2] , \Sum[4][1] ,
         \Sum[4][0] , \Sum[3][31] , \Sum[3][30] , \Sum[3][29] , \Sum[3][28] ,
         \Sum[3][27] , \Sum[3][26] , \Sum[3][25] , \Sum[3][24] , \Sum[3][23] ,
         \Sum[3][22] , \Sum[3][21] , \Sum[3][20] , \Sum[3][19] , \Sum[3][18] ,
         \Sum[3][17] , \Sum[3][16] , \Sum[3][15] , \Sum[3][14] , \Sum[3][13] ,
         \Sum[3][12] , \Sum[3][11] , \Sum[3][10] , \Sum[3][9] , \Sum[3][8] ,
         \Sum[3][7] , \Sum[3][6] , \Sum[3][5] , \Sum[3][4] , \Sum[3][3] ,
         \Sum[3][2] , \Sum[3][1] , \Sum[3][0] , \Sum[2][31] , \Sum[2][30] ,
         \Sum[2][29] , \Sum[2][28] , \Sum[2][27] , \Sum[2][26] , \Sum[2][25] ,
         \Sum[2][24] , \Sum[2][23] , \Sum[2][22] , \Sum[2][21] , \Sum[2][20] ,
         \Sum[2][19] , \Sum[2][18] , \Sum[2][17] , \Sum[2][16] , \Sum[2][15] ,
         \Sum[2][14] , \Sum[2][13] , \Sum[2][12] , \Sum[2][11] , \Sum[2][10] ,
         \Sum[2][9] , \Sum[2][8] , \Sum[2][7] , \Sum[2][6] , \Sum[2][5] ,
         \Sum[2][4] , \Sum[2][3] , \Sum[2][2] , \Sum[2][1] , \Sum[2][0] ,
         \Sum[1][31] , \Sum[1][30] , \Sum[1][29] , \Sum[1][28] , \Sum[1][27] ,
         \Sum[1][26] , \Sum[1][25] , \Sum[1][24] , \Sum[1][23] , \Sum[1][22] ,
         \Sum[1][21] , \Sum[1][20] , \Sum[1][19] , \Sum[1][18] , \Sum[1][17] ,
         \Sum[1][16] , \Sum[1][15] , \Sum[1][14] , \Sum[1][13] , \Sum[1][12] ,
         \Sum[1][11] , \Sum[1][10] , \Sum[1][9] , \Sum[1][8] , \Sum[1][7] ,
         \Sum[1][6] , \Sum[1][5] , \Sum[1][4] , \Sum[1][3] , \Sum[1][2] ,
         \Sum[1][1] , \Sum[1][0] , \Addend[7][31] , \Addend[7][30] ,
         \Addend[7][29] , \Addend[7][28] , \Addend[7][27] , \Addend[7][26] ,
         \Addend[7][25] , \Addend[7][24] , \Addend[7][23] , \Addend[7][22] ,
         \Addend[7][21] , \Addend[7][20] , \Addend[7][19] , \Addend[7][18] ,
         \Addend[7][17] , \Addend[7][16] , \Addend[7][15] , \Addend[7][14] ,
         \Addend[7][13] , \Addend[7][12] , \Addend[7][11] , \Addend[7][10] ,
         \Addend[7][9] , \Addend[7][8] , \Addend[7][7] , \Addend[7][6] ,
         \Addend[7][5] , \Addend[7][4] , \Addend[7][3] , \Addend[7][2] ,
         \Addend[7][1] , \Addend[7][0] , \Addend[6][31] , \Addend[6][30] ,
         \Addend[6][29] , \Addend[6][28] , \Addend[6][27] , \Addend[6][26] ,
         \Addend[6][25] , \Addend[6][24] , \Addend[6][23] , \Addend[6][22] ,
         \Addend[6][21] , \Addend[6][20] , \Addend[6][19] , \Addend[6][18] ,
         \Addend[6][17] , \Addend[6][16] , \Addend[6][15] , \Addend[6][14] ,
         \Addend[6][13] , \Addend[6][12] , \Addend[6][11] , \Addend[6][10] ,
         \Addend[6][9] , \Addend[6][8] , \Addend[6][7] , \Addend[6][6] ,
         \Addend[6][5] , \Addend[6][4] , \Addend[6][3] , \Addend[6][2] ,
         \Addend[6][1] , \Addend[6][0] , \Addend[5][31] , \Addend[5][30] ,
         \Addend[5][29] , \Addend[5][28] , \Addend[5][27] , \Addend[5][26] ,
         \Addend[5][25] , \Addend[5][24] , \Addend[5][23] , \Addend[5][22] ,
         \Addend[5][21] , \Addend[5][20] , \Addend[5][19] , \Addend[5][18] ,
         \Addend[5][17] , \Addend[5][16] , \Addend[5][15] , \Addend[5][14] ,
         \Addend[5][13] , \Addend[5][12] , \Addend[5][11] , \Addend[5][10] ,
         \Addend[5][9] , \Addend[5][8] , \Addend[5][7] , \Addend[5][6] ,
         \Addend[5][5] , \Addend[5][4] , \Addend[5][3] , \Addend[5][2] ,
         \Addend[5][1] , \Addend[5][0] , \Addend[4][31] , \Addend[4][30] ,
         \Addend[4][29] , \Addend[4][28] , \Addend[4][27] , \Addend[4][26] ,
         \Addend[4][25] , \Addend[4][24] , \Addend[4][23] , \Addend[4][22] ,
         \Addend[4][21] , \Addend[4][20] , \Addend[4][19] , \Addend[4][18] ,
         \Addend[4][17] , \Addend[4][16] , \Addend[4][15] , \Addend[4][14] ,
         \Addend[4][13] , \Addend[4][12] , \Addend[4][11] , \Addend[4][10] ,
         \Addend[4][9] , \Addend[4][8] , \Addend[4][7] , \Addend[4][6] ,
         \Addend[4][5] , \Addend[4][4] , \Addend[4][3] , \Addend[4][2] ,
         \Addend[4][1] , \Addend[4][0] , \Addend[3][31] , \Addend[3][30] ,
         \Addend[3][29] , \Addend[3][28] , \Addend[3][27] , \Addend[3][26] ,
         \Addend[3][25] , \Addend[3][24] , \Addend[3][23] , \Addend[3][22] ,
         \Addend[3][21] , \Addend[3][20] , \Addend[3][19] , \Addend[3][18] ,
         \Addend[3][17] , \Addend[3][16] , \Addend[3][15] , \Addend[3][14] ,
         \Addend[3][13] , \Addend[3][12] , \Addend[3][11] , \Addend[3][10] ,
         \Addend[3][9] , \Addend[3][8] , \Addend[3][7] , \Addend[3][6] ,
         \Addend[3][5] , \Addend[3][4] , \Addend[3][3] , \Addend[3][2] ,
         \Addend[3][1] , \Addend[3][0] , \Addend[2][31] , \Addend[2][30] ,
         \Addend[2][29] , \Addend[2][28] , \Addend[2][27] , \Addend[2][26] ,
         \Addend[2][25] , \Addend[2][24] , \Addend[2][23] , \Addend[2][22] ,
         \Addend[2][21] , \Addend[2][20] , \Addend[2][19] , \Addend[2][18] ,
         \Addend[2][17] , \Addend[2][16] , \Addend[2][15] , \Addend[2][14] ,
         \Addend[2][13] , \Addend[2][12] , \Addend[2][11] , \Addend[2][10] ,
         \Addend[2][9] , \Addend[2][8] , \Addend[2][7] , \Addend[2][6] ,
         \Addend[2][5] , \Addend[2][4] , \Addend[2][3] , \Addend[2][2] ,
         \Addend[2][1] , \Addend[2][0] , \Addend[1][31] , \Addend[1][30] ,
         \Addend[1][29] , \Addend[1][28] , \Addend[1][27] , \Addend[1][26] ,
         \Addend[1][25] , \Addend[1][24] , \Addend[1][23] , \Addend[1][22] ,
         \Addend[1][21] , \Addend[1][20] , \Addend[1][19] , \Addend[1][18] ,
         \Addend[1][17] , \Addend[1][16] , \Addend[1][15] , \Addend[1][14] ,
         \Addend[1][13] , \Addend[1][12] , \Addend[1][11] , \Addend[1][10] ,
         \Addend[1][9] , \Addend[1][8] , \Addend[1][7] , \Addend[1][6] ,
         \Addend[1][5] , \Addend[1][4] , \Addend[1][3] , \Addend[1][2] ,
         \Addend[1][1] , \Addend[1][0] , n43, n45, n56, n61, n62, n64, n65,
         n67, n70, n78, n79, n80, n84, n86, n90, n91, n94, n95, n99, n129,
         n146, n158, n160, n163, n168, n172, n174, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20;
  assign n43 = A[7];
  assign n45 = A[1];
  assign n70 = A[3];
  assign n79 = A[4];
  assign n86 = A[6];
  assign n90 = A[0];
  assign n94 = A[5];
  assign n95 = A[8];
  assign n129 = A[15];
  assign n146 = A[2];
  assign n158 = A[9];
  assign n160 = A[10];
  assign n163 = A[11];
  assign n168 = A[12];
  assign n172 = A[13];
  assign n174 = A[14];

  Boothencoder_0 En0_0 ( .B({n286, B[0], 1'b0}), .S({\Sel[0][2] , n99, 
        \Sel[0][0] }) );
  mux51_generic_N32_0 Mux0_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n308, n311, n308, n313, n311, n308, n310, n308, n308, n311, 
        n310, n311, n311, n311, n313, n309, n129, n174, n220, n168, n342, n340, 
        n231, n272, n43, n248, n336, n334, n224, n329, n45, n326}), .C({n297, 
        n295, n297, n297, n297, n298, n297, n297, n296, n295, n298, n297, n299, 
        n295, n299, n299, n56, n279, n78, n280, n227, n65, n382, n212, n64, 
        n262, n84, n223, n264, n91, n61, n325}), .D({n306, n307, n310, n310, 
        n313, n310, n307, n313, n311, n307, n313, n306, n307, n313, n310, n314, 
        n174, n220, n168, n342, n340, n231, n272, n43, n247, n336, n334, n224, 
        n329, n45, n218, 1'b0}), .E({n295, n296, n296, n295, n295, n295, n297, 
        n296, n296, n295, n296, n295, n298, n297, n293, n56, n279, n78, n280, 
        n227, n269, n382, n212, n278, n262, n216, n223, n264, n91, n61, n326, 
        1'b0}), .S({\Sel[0][2] , n99, \Sel[0][0] }), .Y({\Sum[1][31] , 
        \Sum[1][30] , \Sum[1][29] , \Sum[1][28] , \Sum[1][27] , \Sum[1][26] , 
        \Sum[1][25] , \Sum[1][24] , \Sum[1][23] , \Sum[1][22] , \Sum[1][21] , 
        \Sum[1][20] , \Sum[1][19] , \Sum[1][18] , \Sum[1][17] , \Sum[1][16] , 
        \Sum[1][15] , \Sum[1][14] , \Sum[1][13] , \Sum[1][12] , \Sum[1][11] , 
        \Sum[1][10] , \Sum[1][9] , \Sum[1][8] , \Sum[1][7] , \Sum[1][6] , 
        \Sum[1][5] , \Sum[1][4] , \Sum[1][3] , \Sum[1][2] , \Sum[1][1] , 
        \Sum[1][0] }) );
  Boothencoder_7 Eni_1 ( .B(B[3:1]), .S({\Sel[1][2] , \Sel[1][1] , \Sel[1][0] }) );
  mux51_generic_N32_7 Muxi_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n311, n312, n312, n312, n310, n313, n311, n311, n310, n310, 
        n310, n313, n310, n311, n312, n174, n220, n168, n343, n340, n231, n272, 
        n43, n248, n336, n334, n224, n329, n45, n219, 1'b0, 1'b0}), .C({n296, 
        n297, n298, n296, n296, n296, n295, n297, n297, n296, n296, n295, n297, 
        n296, n383, n279, n78, n280, n227, n270, n382, n213, n278, n263, n215, 
        n229, n264, n91, n61, n325, 1'b0, 1'b0}), .D({n307, n308, n307, n307, 
        n307, n308, n307, n308, n308, n313, n308, n313, n310, n308, n174, n172, 
        n168, n342, n340, n231, n272, n43, n247, n336, n334, n224, n329, n45, 
        n324, 1'b0, 1'b0, 1'b0}), .E({n297, n295, n294, n294, n294, n294, n294, 
        n294, n294, n294, n294, n293, n294, n383, n279, n78, n280, n227, n270, 
        n382, n214, n208, n263, n216, n229, n264, n91, n285, n324, 1'b0, 1'b0, 
        1'b0}), .S({\Sel[1][2] , \Sel[1][1] , \Sel[1][0] }), .Y({
        \Addend[1][31] , \Addend[1][30] , \Addend[1][29] , \Addend[1][28] , 
        \Addend[1][27] , \Addend[1][26] , \Addend[1][25] , \Addend[1][24] , 
        \Addend[1][23] , \Addend[1][22] , \Addend[1][21] , \Addend[1][20] , 
        \Addend[1][19] , \Addend[1][18] , \Addend[1][17] , \Addend[1][16] , 
        \Addend[1][15] , \Addend[1][14] , \Addend[1][13] , \Addend[1][12] , 
        \Addend[1][11] , \Addend[1][10] , \Addend[1][9] , \Addend[1][8] , 
        \Addend[1][7] , \Addend[1][6] , \Addend[1][5] , \Addend[1][4] , 
        \Addend[1][3] , \Addend[1][2] , \Addend[1][1] , \Addend[1][0] }) );
  p4adder_N32_7 Addi_1 ( .A({\Addend[1][31] , \Addend[1][30] , \Addend[1][29] , 
        \Addend[1][28] , \Addend[1][27] , \Addend[1][26] , \Addend[1][25] , 
        \Addend[1][24] , \Addend[1][23] , \Addend[1][22] , \Addend[1][21] , 
        \Addend[1][20] , \Addend[1][19] , \Addend[1][18] , \Addend[1][17] , 
        \Addend[1][16] , \Addend[1][15] , \Addend[1][14] , \Addend[1][13] , 
        \Addend[1][12] , \Addend[1][11] , \Addend[1][10] , \Addend[1][9] , 
        n210, \Addend[1][7] , \Addend[1][6] , \Addend[1][5] , \Addend[1][4] , 
        \Addend[1][3] , \Addend[1][2] , \Addend[1][1] , \Addend[1][0] }), .B({
        \Sum[1][31] , \Sum[1][30] , \Sum[1][29] , \Sum[1][28] , \Sum[1][27] , 
        \Sum[1][26] , \Sum[1][25] , \Sum[1][24] , \Sum[1][23] , \Sum[1][22] , 
        \Sum[1][21] , \Sum[1][20] , \Sum[1][19] , \Sum[1][18] , \Sum[1][17] , 
        \Sum[1][16] , \Sum[1][15] , \Sum[1][14] , \Sum[1][13] , \Sum[1][12] , 
        \Sum[1][11] , \Sum[1][10] , \Sum[1][9] , \Sum[1][8] , \Sum[1][7] , 
        \Sum[1][6] , \Sum[1][5] , \Sum[1][4] , \Sum[1][3] , \Sum[1][2] , 
        \Sum[1][1] , \Sum[1][0] }), .Cin(1'b0), .S({\Sum[2][31] , \Sum[2][30] , 
        \Sum[2][29] , \Sum[2][28] , \Sum[2][27] , \Sum[2][26] , \Sum[2][25] , 
        \Sum[2][24] , \Sum[2][23] , \Sum[2][22] , \Sum[2][21] , \Sum[2][20] , 
        \Sum[2][19] , \Sum[2][18] , \Sum[2][17] , \Sum[2][16] , \Sum[2][15] , 
        \Sum[2][14] , \Sum[2][13] , \Sum[2][12] , \Sum[2][11] , \Sum[2][10] , 
        \Sum[2][9] , \Sum[2][8] , \Sum[2][7] , \Sum[2][6] , \Sum[2][5] , 
        \Sum[2][4] , \Sum[2][3] , \Sum[2][2] , \Sum[2][1] , \Sum[2][0] }) );
  Boothencoder_6 Eni_2 ( .B({B[5:4], n221}), .S({\Sel[2][2] , \Sel[2][1] , 
        \Sel[2][0] }) );
  mux51_generic_N32_6 Muxi_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n310, n313, n310, n312, n310, n310, n313, n311, n310, n310, 
        n311, n311, n311, n174, n220, n168, n342, n340, n231, n272, n43, n247, 
        n336, n334, n224, n329, n45, n218, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n294, 
        n293, n293, n293, n293, n293, n293, n293, n293, n293, n293, n293, n244, 
        n279, n78, n280, n275, n270, n382, n214, n226, n263, n215, n246, n253, 
        n256, n285, n325, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n312, n309, n312, n310, 
        n311, n312, n310, n310, n310, n313, n313, n313, n174, n172, n168, n342, 
        n340, n231, n272, n43, n248, n336, n334, n224, n329, n45, n219, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .E({n292, n292, n292, n292, n292, n292, n292, 
        n292, n292, n292, n292, n245, n279, n78, n280, n275, n270, n382, n213, 
        n208, n263, n216, n246, n253, n91, n285, n326, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S({\Sel[2][2] , \Sel[2][1] , \Sel[2][0] }), .Y({
        \Addend[2][31] , \Addend[2][30] , \Addend[2][29] , \Addend[2][28] , 
        \Addend[2][27] , \Addend[2][26] , \Addend[2][25] , \Addend[2][24] , 
        \Addend[2][23] , \Addend[2][22] , \Addend[2][21] , \Addend[2][20] , 
        \Addend[2][19] , \Addend[2][18] , \Addend[2][17] , \Addend[2][16] , 
        \Addend[2][15] , \Addend[2][14] , \Addend[2][13] , \Addend[2][12] , 
        \Addend[2][11] , \Addend[2][10] , \Addend[2][9] , \Addend[2][8] , 
        \Addend[2][7] , \Addend[2][6] , \Addend[2][5] , \Addend[2][4] , 
        \Addend[2][3] , \Addend[2][2] , \Addend[2][1] , \Addend[2][0] }) );
  p4adder_N32_6 Addi_2 ( .A({\Addend[2][31] , \Addend[2][30] , \Addend[2][29] , 
        \Addend[2][28] , \Addend[2][27] , \Addend[2][26] , \Addend[2][25] , 
        \Addend[2][24] , \Addend[2][23] , \Addend[2][22] , \Addend[2][21] , 
        \Addend[2][20] , \Addend[2][19] , \Addend[2][18] , \Addend[2][17] , 
        \Addend[2][16] , \Addend[2][15] , \Addend[2][14] , \Addend[2][13] , 
        \Addend[2][12] , \Addend[2][11] , \Addend[2][10] , \Addend[2][9] , 
        \Addend[2][8] , \Addend[2][7] , \Addend[2][6] , \Addend[2][5] , 
        \Addend[2][4] , \Addend[2][3] , \Addend[2][2] , \Addend[2][1] , 
        \Addend[2][0] }), .B({\Sum[2][31] , \Sum[2][30] , \Sum[2][29] , 
        \Sum[2][28] , \Sum[2][27] , \Sum[2][26] , \Sum[2][25] , \Sum[2][24] , 
        \Sum[2][23] , \Sum[2][22] , \Sum[2][21] , \Sum[2][20] , \Sum[2][19] , 
        \Sum[2][18] , \Sum[2][17] , \Sum[2][16] , \Sum[2][15] , \Sum[2][14] , 
        \Sum[2][13] , \Sum[2][12] , \Sum[2][11] , \Sum[2][10] , \Sum[2][9] , 
        \Sum[2][8] , \Sum[2][7] , \Sum[2][6] , \Sum[2][5] , \Sum[2][4] , 
        \Sum[2][3] , \Sum[2][2] , \Sum[2][1] , \Sum[2][0] }), .Cin(1'b0), .S({
        \Sum[3][31] , \Sum[3][30] , \Sum[3][29] , \Sum[3][28] , \Sum[3][27] , 
        \Sum[3][26] , \Sum[3][25] , \Sum[3][24] , \Sum[3][23] , \Sum[3][22] , 
        \Sum[3][21] , \Sum[3][20] , \Sum[3][19] , \Sum[3][18] , \Sum[3][17] , 
        \Sum[3][16] , \Sum[3][15] , \Sum[3][14] , \Sum[3][13] , \Sum[3][12] , 
        \Sum[3][11] , \Sum[3][10] , \Sum[3][9] , \Sum[3][8] , \Sum[3][7] , 
        \Sum[3][6] , \Sum[3][5] , \Sum[3][4] , \Sum[3][3] , \Sum[3][2] , 
        \Sum[3][1] , \Sum[3][0] }) );
  Boothencoder_5 Eni_3 ( .B(B[7:5]), .S({\Sel[3][2] , \Sel[3][1] , \Sel[3][0] }) );
  mux51_generic_N32_5 Muxi_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n310, n311, n313, n309, n309, n309, n312, n311, n313, n310, 
        n310, n174, n220, n168, n342, n340, n231, n272, n43, n248, n336, n334, 
        n224, n329, n45, n219, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n290, 
        n291, n291, n291, n291, n291, n290, n291, n290, n291, n244, n279, n78, 
        n280, n275, n270, n382, n213, n208, n263, n215, n246, n253, n256, n285, 
        n325, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n313, n309, n310, n310, 
        n310, n313, n310, n313, n310, n310, n174, n172, n168, n342, n340, n231, 
        n272, n43, n247, n336, n334, n224, n329, n207, n326, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .E({n290, n289, n290, n290, n290, n290, n290, 
        n290, n289, n245, n279, n78, n280, n275, n270, n382, n214, n226, n263, 
        n216, n246, n253, n256, n285, n218, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S({\Sel[3][2] , \Sel[3][1] , \Sel[3][0] }), .Y({
        \Addend[3][31] , \Addend[3][30] , \Addend[3][29] , \Addend[3][28] , 
        \Addend[3][27] , \Addend[3][26] , \Addend[3][25] , \Addend[3][24] , 
        \Addend[3][23] , \Addend[3][22] , \Addend[3][21] , \Addend[3][20] , 
        \Addend[3][19] , \Addend[3][18] , \Addend[3][17] , \Addend[3][16] , 
        \Addend[3][15] , \Addend[3][14] , \Addend[3][13] , \Addend[3][12] , 
        \Addend[3][11] , \Addend[3][10] , \Addend[3][9] , \Addend[3][8] , 
        \Addend[3][7] , \Addend[3][6] , \Addend[3][5] , \Addend[3][4] , 
        \Addend[3][3] , \Addend[3][2] , \Addend[3][1] , \Addend[3][0] }) );
  p4adder_N32_5 Addi_3 ( .A({\Addend[3][31] , \Addend[3][30] , \Addend[3][29] , 
        \Addend[3][28] , \Addend[3][27] , \Addend[3][26] , \Addend[3][25] , 
        \Addend[3][24] , \Addend[3][23] , \Addend[3][22] , \Addend[3][21] , 
        \Addend[3][20] , \Addend[3][19] , \Addend[3][18] , \Addend[3][17] , 
        \Addend[3][16] , \Addend[3][15] , \Addend[3][14] , \Addend[3][13] , 
        \Addend[3][12] , \Addend[3][11] , \Addend[3][10] , \Addend[3][9] , 
        \Addend[3][8] , \Addend[3][7] , \Addend[3][6] , \Addend[3][5] , 
        \Addend[3][4] , \Addend[3][3] , \Addend[3][2] , \Addend[3][1] , 
        \Addend[3][0] }), .B({\Sum[3][31] , \Sum[3][30] , \Sum[3][29] , 
        \Sum[3][28] , \Sum[3][27] , \Sum[3][26] , \Sum[3][25] , \Sum[3][24] , 
        \Sum[3][23] , \Sum[3][22] , \Sum[3][21] , \Sum[3][20] , \Sum[3][19] , 
        \Sum[3][18] , \Sum[3][17] , \Sum[3][16] , \Sum[3][15] , \Sum[3][14] , 
        \Sum[3][13] , \Sum[3][12] , \Sum[3][11] , \Sum[3][10] , \Sum[3][9] , 
        \Sum[3][8] , \Sum[3][7] , \Sum[3][6] , \Sum[3][5] , \Sum[3][4] , 
        \Sum[3][3] , \Sum[3][2] , \Sum[3][1] , \Sum[3][0] }), .Cin(1'b0), .S({
        \Sum[4][31] , \Sum[4][30] , \Sum[4][29] , \Sum[4][28] , \Sum[4][27] , 
        \Sum[4][26] , \Sum[4][25] , \Sum[4][24] , \Sum[4][23] , \Sum[4][22] , 
        \Sum[4][21] , \Sum[4][20] , \Sum[4][19] , \Sum[4][18] , \Sum[4][17] , 
        \Sum[4][16] , \Sum[4][15] , \Sum[4][14] , \Sum[4][13] , \Sum[4][12] , 
        \Sum[4][11] , \Sum[4][10] , \Sum[4][9] , \Sum[4][8] , \Sum[4][7] , 
        \Sum[4][6] , \Sum[4][5] , \Sum[4][4] , \Sum[4][3] , \Sum[4][2] , 
        \Sum[4][1] , \Sum[4][0] }) );
  Boothencoder_4 Eni_4 ( .B(B[9:7]), .S({\Sel[4][2] , \Sel[4][1] , \Sel[4][0] }) );
  mux51_generic_N32_4 Muxi_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n309, n309, n309, n312, n311, n309, n312, n312, n310, n174, 
        n172, n168, n342, n340, n231, n272, n43, n248, n336, n334, n224, n329, 
        n207, n219, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n290, 
        n289, n290, n289, n289, n289, n289, n289, n245, n279, n78, n276, n275, 
        n270, n382, n213, n226, n263, n215, n246, n253, n256, n285, n326, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n314, n314, n314, n314, 
        n314, n314, n314, n314, n174, n220, n168, n342, n340, n231, n272, n43, 
        n247, n336, n334, n224, n329, n207, n218, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .E({\MinusAExt2[4][31] , \MinusAExt2[4][30] , 
        \MinusAExt2[4][29] , \MinusAExt2[4][28] , \MinusAExt2[4][27] , 
        \MinusAExt2[4][26] , \MinusAExt2[4][25] , \MinusAExt2[4][24] , 
        \MinusAExt2[4][23] , \MinusAExt2[4][22] , \MinusAExt2[4][21] , 
        \MinusAExt2[4][20] , \MinusAExt2[4][19] , \MinusAExt2[4][18] , 
        \MinusAExt2[4][17] , \MinusAExt2[4][16] , \MinusAExt2[4][15] , 
        \MinusAExt2[4][14] , \MinusAExt2[4][13] , \MinusAExt2[4][12] , 
        \MinusAExt2[4][11] , \MinusAExt2[4][10] , \MinusAExt2[4][9] , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S({\Sel[4][2] , 
        \Sel[4][1] , \Sel[4][0] }), .Y({\Addend[4][31] , \Addend[4][30] , 
        \Addend[4][29] , \Addend[4][28] , \Addend[4][27] , \Addend[4][26] , 
        \Addend[4][25] , \Addend[4][24] , \Addend[4][23] , \Addend[4][22] , 
        \Addend[4][21] , \Addend[4][20] , \Addend[4][19] , \Addend[4][18] , 
        \Addend[4][17] , \Addend[4][16] , \Addend[4][15] , \Addend[4][14] , 
        \Addend[4][13] , \Addend[4][12] , \Addend[4][11] , \Addend[4][10] , 
        \Addend[4][9] , \Addend[4][8] , \Addend[4][7] , \Addend[4][6] , 
        \Addend[4][5] , \Addend[4][4] , \Addend[4][3] , \Addend[4][2] , 
        \Addend[4][1] , \Addend[4][0] }) );
  p4adder_N32_4 Addi_4 ( .A({\Addend[4][31] , \Addend[4][30] , \Addend[4][29] , 
        \Addend[4][28] , \Addend[4][27] , \Addend[4][26] , \Addend[4][25] , 
        \Addend[4][24] , \Addend[4][23] , \Addend[4][22] , \Addend[4][21] , 
        \Addend[4][20] , \Addend[4][19] , \Addend[4][18] , \Addend[4][17] , 
        \Addend[4][16] , \Addend[4][15] , \Addend[4][14] , \Addend[4][13] , 
        \Addend[4][12] , \Addend[4][11] , \Addend[4][10] , \Addend[4][9] , 
        \Addend[4][8] , \Addend[4][7] , \Addend[4][6] , \Addend[4][5] , 
        \Addend[4][4] , \Addend[4][3] , \Addend[4][2] , \Addend[4][1] , 
        \Addend[4][0] }), .B({\Sum[4][31] , \Sum[4][30] , \Sum[4][29] , 
        \Sum[4][28] , \Sum[4][27] , \Sum[4][26] , \Sum[4][25] , \Sum[4][24] , 
        \Sum[4][23] , \Sum[4][22] , \Sum[4][21] , \Sum[4][20] , \Sum[4][19] , 
        \Sum[4][18] , \Sum[4][17] , \Sum[4][16] , \Sum[4][15] , \Sum[4][14] , 
        \Sum[4][13] , \Sum[4][12] , \Sum[4][11] , \Sum[4][10] , \Sum[4][9] , 
        \Sum[4][8] , \Sum[4][7] , \Sum[4][6] , \Sum[4][5] , \Sum[4][4] , 
        \Sum[4][3] , \Sum[4][2] , \Sum[4][1] , \Sum[4][0] }), .Cin(1'b0), .S({
        \Sum[5][31] , \Sum[5][30] , \Sum[5][29] , \Sum[5][28] , \Sum[5][27] , 
        \Sum[5][26] , \Sum[5][25] , \Sum[5][24] , \Sum[5][23] , \Sum[5][22] , 
        \Sum[5][21] , \Sum[5][20] , \Sum[5][19] , \Sum[5][18] , \Sum[5][17] , 
        \Sum[5][16] , \Sum[5][15] , \Sum[5][14] , \Sum[5][13] , \Sum[5][12] , 
        \Sum[5][11] , \Sum[5][10] , \Sum[5][9] , \Sum[5][8] , \Sum[5][7] , 
        \Sum[5][6] , \Sum[5][5] , \Sum[5][4] , \Sum[5][3] , \Sum[5][2] , 
        \Sum[5][1] , \Sum[5][0] }) );
  Boothencoder_3 Eni_5 ( .B(B[11:9]), .S({\Sel[5][2] , \Sel[5][1] , 
        \Sel[5][0] }) );
  mux51_generic_N32_3 Muxi_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n310, n311, n314, n313, n308, n309, n311, n174, n220, n168, 
        n342, n340, n231, n272, n43, n248, n336, n334, n224, n329, n207, n326, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({
        \MinusAExt1[5][31] , \MinusAExt1[5][30] , \MinusAExt1[5][29] , 
        \MinusAExt1[5][28] , \MinusAExt1[5][27] , \MinusAExt1[5][26] , 
        \MinusAExt1[5][25] , \MinusAExt1[5][24] , \MinusAExt1[5][23] , 
        \MinusAExt1[5][22] , \MinusAExt1[5][21] , \MinusAExt1[5][20] , 
        \MinusAExt1[5][19] , \MinusAExt1[5][18] , \MinusAExt1[5][17] , 
        \MinusAExt1[5][16] , \MinusAExt1[5][15] , \MinusAExt1[5][14] , 
        \MinusAExt1[5][13] , \MinusAExt1[5][12] , \MinusAExt1[5][11] , 
        \MinusAExt1[5][10] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .D({n309, n310, n310, n312, n307, n310, n174, n172, n168, 
        n342, n340, n231, n272, n43, n247, n336, n334, n224, n329, n207, n325, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .E({n289, n289, n289, n289, n298, n244, n279, n78, n233, n275, n270, 
        n242, n214, n208, n263, n216, n246, n253, n256, n285, n219, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S({
        \Sel[5][2] , \Sel[5][1] , \Sel[5][0] }), .Y({\Addend[5][31] , 
        \Addend[5][30] , \Addend[5][29] , \Addend[5][28] , \Addend[5][27] , 
        \Addend[5][26] , \Addend[5][25] , \Addend[5][24] , \Addend[5][23] , 
        \Addend[5][22] , \Addend[5][21] , \Addend[5][20] , \Addend[5][19] , 
        \Addend[5][18] , \Addend[5][17] , \Addend[5][16] , \Addend[5][15] , 
        \Addend[5][14] , \Addend[5][13] , \Addend[5][12] , \Addend[5][11] , 
        \Addend[5][10] , \Addend[5][9] , \Addend[5][8] , \Addend[5][7] , 
        \Addend[5][6] , \Addend[5][5] , \Addend[5][4] , \Addend[5][3] , 
        \Addend[5][2] , \Addend[5][1] , \Addend[5][0] }) );
  p4adder_N32_3 Addi_5 ( .A({\Addend[5][31] , \Addend[5][30] , \Addend[5][29] , 
        \Addend[5][28] , \Addend[5][27] , \Addend[5][26] , \Addend[5][25] , 
        \Addend[5][24] , \Addend[5][23] , \Addend[5][22] , \Addend[5][21] , 
        \Addend[5][20] , \Addend[5][19] , \Addend[5][18] , \Addend[5][17] , 
        \Addend[5][16] , \Addend[5][15] , \Addend[5][14] , \Addend[5][13] , 
        \Addend[5][12] , \Addend[5][11] , \Addend[5][10] , \Addend[5][9] , 
        \Addend[5][8] , \Addend[5][7] , \Addend[5][6] , \Addend[5][5] , 
        \Addend[5][4] , \Addend[5][3] , \Addend[5][2] , \Addend[5][1] , 
        \Addend[5][0] }), .B({\Sum[5][31] , \Sum[5][30] , \Sum[5][29] , 
        \Sum[5][28] , \Sum[5][27] , \Sum[5][26] , \Sum[5][25] , \Sum[5][24] , 
        \Sum[5][23] , \Sum[5][22] , \Sum[5][21] , \Sum[5][20] , \Sum[5][19] , 
        \Sum[5][18] , \Sum[5][17] , \Sum[5][16] , \Sum[5][15] , \Sum[5][14] , 
        \Sum[5][13] , \Sum[5][12] , \Sum[5][11] , \Sum[5][10] , \Sum[5][9] , 
        \Sum[5][8] , \Sum[5][7] , \Sum[5][6] , \Sum[5][5] , \Sum[5][4] , 
        \Sum[5][3] , \Sum[5][2] , \Sum[5][1] , \Sum[5][0] }), .Cin(1'b0), .S({
        \Sum[6][31] , \Sum[6][30] , \Sum[6][29] , \Sum[6][28] , \Sum[6][27] , 
        \Sum[6][26] , \Sum[6][25] , \Sum[6][24] , \Sum[6][23] , \Sum[6][22] , 
        \Sum[6][21] , \Sum[6][20] , \Sum[6][19] , \Sum[6][18] , \Sum[6][17] , 
        \Sum[6][16] , \Sum[6][15] , \Sum[6][14] , \Sum[6][13] , \Sum[6][12] , 
        \Sum[6][11] , \Sum[6][10] , \Sum[6][9] , \Sum[6][8] , \Sum[6][7] , 
        \Sum[6][6] , \Sum[6][5] , \Sum[6][4] , \Sum[6][3] , \Sum[6][2] , 
        \Sum[6][1] , \Sum[6][0] }) );
  Boothencoder_2 Eni_6 ( .B(B[13:11]), .S({\Sel[6][2] , \Sel[6][1] , 
        \Sel[6][0] }) );
  mux51_generic_N32_2 Muxi_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n307, n307, n306, n306, n312, n174, n172, n168, n342, n340, 
        n231, n272, n43, n248, n336, n334, n224, n329, n207, n325, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n291, 
        n291, n292, n291, n244, n279, n78, n233, n275, n270, n382, n230, n281, 
        n263, n236, n246, n253, n256, n285, n218, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n306, n306, n306, n306, 
        n174, n220, n168, n342, n340, n231, n272, n43, n247, n336, n334, n224, 
        n329, n207, n219, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .E({n297, n295, n296, n245, n279, n78, n233, 
        n275, n270, n242, n214, n281, n263, n236, n246, n253, n256, n285, n218, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S({\Sel[6][2] , \Sel[6][1] , \Sel[6][0] }), .Y({
        \Addend[6][31] , \Addend[6][30] , \Addend[6][29] , \Addend[6][28] , 
        \Addend[6][27] , \Addend[6][26] , \Addend[6][25] , \Addend[6][24] , 
        \Addend[6][23] , \Addend[6][22] , \Addend[6][21] , \Addend[6][20] , 
        \Addend[6][19] , \Addend[6][18] , \Addend[6][17] , \Addend[6][16] , 
        \Addend[6][15] , \Addend[6][14] , \Addend[6][13] , \Addend[6][12] , 
        \Addend[6][11] , \Addend[6][10] , \Addend[6][9] , \Addend[6][8] , 
        \Addend[6][7] , \Addend[6][6] , \Addend[6][5] , \Addend[6][4] , 
        \Addend[6][3] , \Addend[6][2] , \Addend[6][1] , \Addend[6][0] }) );
  p4adder_N32_2 Addi_6 ( .A({\Addend[6][31] , \Addend[6][30] , \Addend[6][29] , 
        \Addend[6][28] , \Addend[6][27] , \Addend[6][26] , \Addend[6][25] , 
        \Addend[6][24] , \Addend[6][23] , \Addend[6][22] , \Addend[6][21] , 
        \Addend[6][20] , \Addend[6][19] , \Addend[6][18] , \Addend[6][17] , 
        \Addend[6][16] , \Addend[6][15] , \Addend[6][14] , \Addend[6][13] , 
        \Addend[6][12] , \Addend[6][11] , \Addend[6][10] , \Addend[6][9] , 
        \Addend[6][8] , \Addend[6][7] , \Addend[6][6] , \Addend[6][5] , 
        \Addend[6][4] , \Addend[6][3] , \Addend[6][2] , \Addend[6][1] , 
        \Addend[6][0] }), .B({\Sum[6][31] , \Sum[6][30] , \Sum[6][29] , 
        \Sum[6][28] , \Sum[6][27] , \Sum[6][26] , \Sum[6][25] , \Sum[6][24] , 
        \Sum[6][23] , \Sum[6][22] , \Sum[6][21] , \Sum[6][20] , \Sum[6][19] , 
        \Sum[6][18] , \Sum[6][17] , \Sum[6][16] , \Sum[6][15] , \Sum[6][14] , 
        \Sum[6][13] , \Sum[6][12] , \Sum[6][11] , \Sum[6][10] , \Sum[6][9] , 
        \Sum[6][8] , \Sum[6][7] , \Sum[6][6] , \Sum[6][5] , \Sum[6][4] , 
        \Sum[6][3] , \Sum[6][2] , \Sum[6][1] , \Sum[6][0] }), .Cin(1'b0), .S({
        \Sum[7][31] , \Sum[7][30] , \Sum[7][29] , \Sum[7][28] , \Sum[7][27] , 
        \Sum[7][26] , \Sum[7][25] , \Sum[7][24] , \Sum[7][23] , \Sum[7][22] , 
        \Sum[7][21] , \Sum[7][20] , \Sum[7][19] , \Sum[7][18] , \Sum[7][17] , 
        \Sum[7][16] , \Sum[7][15] , \Sum[7][14] , \Sum[7][13] , \Sum[7][12] , 
        \Sum[7][11] , \Sum[7][10] , \Sum[7][9] , \Sum[7][8] , \Sum[7][7] , 
        \Sum[7][6] , \Sum[7][5] , \Sum[7][4] , \Sum[7][3] , \Sum[7][2] , 
        \Sum[7][1] , \Sum[7][0] }) );
  Boothencoder_1 Eni_7 ( .B(B[15:13]), .S({\Sel[7][2] , \Sel[7][1] , 
        \Sel[7][0] }) );
  mux51_generic_N32_1 Muxi_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .B({n306, n306, n312, n174, n220, n168, n342, n340, n231, n272, 
        n43, n247, n336, n334, n224, n329, n207, n238, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n291, 
        n291, n244, n279, n78, n280, n275, n270, n242, n230, n281, n263, n236, 
        n246, n253, n256, n285, n219, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n306, n306, n174, n172, 
        n168, n342, n340, n231, n272, n43, n248, n336, n334, n224, n329, n207, 
        n218, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .E({n298, n245, n279, n78, n276, n275, n270, 
        n242, n230, n281, n263, n236, n246, n253, n256, n285, n325, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S({\Sel[7][2] , \Sel[7][1] , \Sel[7][0] }), .Y({
        \Addend[7][31] , \Addend[7][30] , \Addend[7][29] , \Addend[7][28] , 
        \Addend[7][27] , \Addend[7][26] , \Addend[7][25] , \Addend[7][24] , 
        \Addend[7][23] , \Addend[7][22] , \Addend[7][21] , \Addend[7][20] , 
        \Addend[7][19] , \Addend[7][18] , \Addend[7][17] , \Addend[7][16] , 
        \Addend[7][15] , \Addend[7][14] , \Addend[7][13] , \Addend[7][12] , 
        \Addend[7][11] , \Addend[7][10] , \Addend[7][9] , \Addend[7][8] , 
        \Addend[7][7] , \Addend[7][6] , \Addend[7][5] , \Addend[7][4] , 
        \Addend[7][3] , \Addend[7][2] , \Addend[7][1] , \Addend[7][0] }) );
  p4adder_N32_1 Addi_7 ( .A({\Addend[7][31] , \Addend[7][30] , \Addend[7][29] , 
        \Addend[7][28] , \Addend[7][27] , \Addend[7][26] , \Addend[7][25] , 
        \Addend[7][24] , \Addend[7][23] , \Addend[7][22] , \Addend[7][21] , 
        \Addend[7][20] , \Addend[7][19] , \Addend[7][18] , \Addend[7][17] , 
        \Addend[7][16] , \Addend[7][15] , \Addend[7][14] , \Addend[7][13] , 
        \Addend[7][12] , \Addend[7][11] , \Addend[7][10] , \Addend[7][9] , 
        \Addend[7][8] , \Addend[7][7] , \Addend[7][6] , \Addend[7][5] , 
        \Addend[7][4] , \Addend[7][3] , \Addend[7][2] , \Addend[7][1] , 
        \Addend[7][0] }), .B({\Sum[7][31] , \Sum[7][30] , \Sum[7][29] , 
        \Sum[7][28] , \Sum[7][27] , \Sum[7][26] , \Sum[7][25] , \Sum[7][24] , 
        \Sum[7][23] , \Sum[7][22] , \Sum[7][21] , \Sum[7][20] , \Sum[7][19] , 
        \Sum[7][18] , \Sum[7][17] , \Sum[7][16] , \Sum[7][15] , \Sum[7][14] , 
        \Sum[7][13] , \Sum[7][12] , \Sum[7][11] , \Sum[7][10] , \Sum[7][9] , 
        \Sum[7][8] , \Sum[7][7] , \Sum[7][6] , \Sum[7][5] , \Sum[7][4] , 
        \Sum[7][3] , \Sum[7][2] , \Sum[7][1] , \Sum[7][0] }), .Cin(1'b0), .S(P) );
  Boothmul_N16_DW01_inc_5 add_74_G6 ( .A({1'b0, n318, n315, n315, n315, n315, 
        n316, n316, n350, n349, n347, n345, n341, n235, n338, n241, n305, n258, 
        n243, n333, n332, n261, n217, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .SUM({SYNOPSYS_UNCONNECTED__0, \MinusAExt1[5][31] , 
        \MinusAExt1[5][30] , \MinusAExt1[5][29] , \MinusAExt1[5][28] , 
        \MinusAExt1[5][27] , \MinusAExt1[5][26] , \MinusAExt1[5][25] , 
        \MinusAExt1[5][24] , \MinusAExt1[5][23] , \MinusAExt1[5][22] , 
        \MinusAExt1[5][21] , \MinusAExt1[5][20] , \MinusAExt1[5][19] , 
        \MinusAExt1[5][18] , \MinusAExt1[5][17] , \MinusAExt1[5][16] , 
        \MinusAExt1[5][15] , \MinusAExt1[5][14] , \MinusAExt1[5][13] , 
        \MinusAExt1[5][12] , \MinusAExt1[5][11] , \MinusAExt1[5][10] , 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10}) );
  Boothmul_N16_DW01_inc_6 add_76_G5 ( .A({1'b0, n318, n316, n316, n317, n317, 
        n317, n317, n318, n350, n349, n347, n345, n341, n235, n338, n241, n304, 
        n258, n243, n333, n332, n261, n217, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1}), .SUM({SYNOPSYS_UNCONNECTED__11, 
        \MinusAExt2[4][31] , \MinusAExt2[4][30] , \MinusAExt2[4][29] , 
        \MinusAExt2[4][28] , \MinusAExt2[4][27] , \MinusAExt2[4][26] , 
        \MinusAExt2[4][25] , \MinusAExt2[4][24] , \MinusAExt2[4][23] , 
        \MinusAExt2[4][22] , \MinusAExt2[4][21] , \MinusAExt2[4][20] , 
        \MinusAExt2[4][19] , \MinusAExt2[4][18] , \MinusAExt2[4][17] , 
        \MinusAExt2[4][16] , \MinusAExt2[4][15] , \MinusAExt2[4][14] , 
        \MinusAExt2[4][13] , \MinusAExt2[4][12] , \MinusAExt2[4][11] , 
        \MinusAExt2[4][10] , \MinusAExt2[4][9] , SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20}) );
  XNOR2_X1 U3 ( .A(n266), .B(n160), .ZN(n65) );
  CLKBUF_X1 U4 ( .A(n45), .Z(n207) );
  INV_X1 U5 ( .A(n352), .ZN(n285) );
  CLKBUF_X1 U6 ( .A(n91), .Z(n256) );
  AND2_X2 U7 ( .A1(n356), .A2(n357), .ZN(n264) );
  INV_X1 U8 ( .A(n277), .ZN(n208) );
  CLKBUF_X3 U9 ( .A(n67), .Z(n263) );
  AND3_X2 U10 ( .A1(n361), .A2(n362), .A3(n268), .ZN(n282) );
  AND2_X1 U11 ( .A1(n348), .A2(n346), .ZN(n209) );
  BUF_X2 U12 ( .A(B[1]), .Z(n286) );
  BUF_X1 U13 ( .A(n80), .Z(n213) );
  BUF_X1 U14 ( .A(n327), .Z(n274) );
  BUF_X2 U15 ( .A(n321), .Z(n319) );
  CLKBUF_X1 U16 ( .A(n65), .Z(n269) );
  CLKBUF_X3 U17 ( .A(n65), .Z(n270) );
  BUF_X1 U18 ( .A(n381), .Z(n288) );
  BUF_X1 U19 ( .A(n381), .Z(n287) );
  BUF_X1 U20 ( .A(n67), .Z(n262) );
  BUF_X2 U21 ( .A(\Addend[1][8] ), .Z(n210) );
  INV_X1 U22 ( .A(n146), .ZN(n211) );
  BUF_X1 U23 ( .A(n80), .Z(n212) );
  BUF_X1 U24 ( .A(n80), .Z(n214) );
  XNOR2_X1 U25 ( .A(n363), .B(n272), .ZN(n80) );
  XNOR2_X1 U26 ( .A(n251), .B(n228), .ZN(n216) );
  XNOR2_X1 U27 ( .A(n251), .B(n228), .ZN(n215) );
  AND3_X2 U28 ( .A1(n243), .A2(n265), .A3(n358), .ZN(n251) );
  XNOR2_X1 U29 ( .A(n251), .B(n228), .ZN(n84) );
  INV_X1 U30 ( .A(n90), .ZN(n217) );
  INV_X1 U31 ( .A(n217), .ZN(n219) );
  INV_X1 U32 ( .A(n217), .ZN(n218) );
  BUF_X2 U33 ( .A(n172), .Z(n220) );
  CLKBUF_X1 U34 ( .A(B[3]), .Z(n221) );
  INV_X1 U35 ( .A(n45), .ZN(n222) );
  XNOR2_X1 U36 ( .A(n357), .B(n243), .ZN(n223) );
  XNOR2_X1 U37 ( .A(n357), .B(n243), .ZN(n229) );
  INV_X2 U38 ( .A(n333), .ZN(n224) );
  OR2_X1 U39 ( .A1(n295), .A2(n378), .ZN(n245) );
  OR2_X1 U40 ( .A1(n295), .A2(n378), .ZN(n244) );
  AND2_X1 U41 ( .A1(n255), .A2(n341), .ZN(n225) );
  AND2_X1 U42 ( .A1(n255), .A2(n341), .ZN(n369) );
  INV_X1 U43 ( .A(n172), .ZN(n349) );
  INV_X1 U44 ( .A(n277), .ZN(n226) );
  AND2_X2 U45 ( .A1(n335), .A2(n331), .ZN(n268) );
  INV_X1 U46 ( .A(n335), .ZN(n334) );
  XNOR2_X1 U47 ( .A(n370), .B(n344), .ZN(n227) );
  CLKBUF_X1 U48 ( .A(n94), .Z(n228) );
  BUF_X2 U49 ( .A(n288), .Z(n293) );
  INV_X1 U50 ( .A(n229), .ZN(n239) );
  BUF_X2 U51 ( .A(n287), .Z(n296) );
  BUF_X1 U52 ( .A(n213), .Z(n230) );
  CLKBUF_X3 U53 ( .A(n158), .Z(n231) );
  NAND2_X1 U54 ( .A1(n225), .A2(n259), .ZN(n232) );
  CLKBUF_X1 U55 ( .A(n280), .Z(n233) );
  INV_X1 U56 ( .A(n86), .ZN(n234) );
  BUF_X1 U57 ( .A(n339), .Z(n235) );
  CLKBUF_X1 U58 ( .A(n215), .Z(n236) );
  INV_X1 U59 ( .A(n326), .ZN(n237) );
  INV_X1 U60 ( .A(n237), .ZN(n238) );
  BUF_X1 U61 ( .A(n327), .Z(n273) );
  INV_X1 U62 ( .A(n354), .ZN(n240) );
  AND2_X1 U63 ( .A1(n222), .A2(n274), .ZN(n265) );
  INV_X1 U64 ( .A(n43), .ZN(n241) );
  CLKBUF_X1 U65 ( .A(n382), .Z(n242) );
  INV_X1 U66 ( .A(n303), .ZN(n301) );
  INV_X1 U67 ( .A(n79), .ZN(n243) );
  INV_X1 U68 ( .A(n79), .ZN(n335) );
  OR2_X1 U69 ( .A1(n299), .A2(n378), .ZN(n383) );
  AND2_X1 U70 ( .A1(n257), .A2(n366), .ZN(n260) );
  INV_X1 U71 ( .A(n239), .ZN(n246) );
  CLKBUF_X3 U72 ( .A(n95), .Z(n272) );
  INV_X1 U193 ( .A(n234), .ZN(n248) );
  INV_X1 U194 ( .A(n234), .ZN(n247) );
  INV_X4 U195 ( .A(n319), .ZN(n310) );
  CLKBUF_X1 U196 ( .A(n95), .Z(n271) );
  NOR2_X1 U197 ( .A1(n249), .A2(n250), .ZN(n255) );
  NAND2_X1 U198 ( .A1(n339), .A2(n267), .ZN(n249) );
  NAND2_X1 U199 ( .A1(n300), .A2(n303), .ZN(n250) );
  INV_X1 U200 ( .A(n264), .ZN(n252) );
  INV_X1 U201 ( .A(n252), .ZN(n253) );
  INV_X1 U202 ( .A(n43), .ZN(n300) );
  AND2_X1 U203 ( .A1(n369), .A2(n282), .ZN(n254) );
  XNOR2_X1 U204 ( .A(n355), .B(n332), .ZN(n91) );
  AND3_X1 U205 ( .A1(n359), .A2(n268), .A3(n265), .ZN(n257) );
  INV_X1 U206 ( .A(n336), .ZN(n258) );
  NAND2_X1 U207 ( .A1(n225), .A2(n259), .ZN(n374) );
  AND2_X1 U208 ( .A1(n282), .A2(n209), .ZN(n259) );
  XNOR2_X2 U209 ( .A(n260), .B(n158), .ZN(n382) );
  INV_X1 U210 ( .A(n337), .ZN(n336) );
  INV_X1 U211 ( .A(n94), .ZN(n337) );
  INV_X1 U212 ( .A(n45), .ZN(n261) );
  XNOR2_X1 U213 ( .A(n364), .B(n305), .ZN(n67) );
  CLKBUF_X1 U214 ( .A(n287), .Z(n298) );
  BUF_X1 U215 ( .A(n288), .Z(n299) );
  BUF_X1 U216 ( .A(n322), .Z(n318) );
  CLKBUF_X1 U217 ( .A(n287), .Z(n292) );
  BUF_X2 U218 ( .A(n288), .Z(n295) );
  BUF_X1 U219 ( .A(n287), .Z(n294) );
  BUF_X2 U220 ( .A(n288), .Z(n297) );
  CLKBUF_X1 U221 ( .A(n287), .Z(n289) );
  CLKBUF_X1 U222 ( .A(n287), .Z(n290) );
  CLKBUF_X1 U223 ( .A(n287), .Z(n291) );
  INV_X1 U224 ( .A(n319), .ZN(n311) );
  INV_X1 U225 ( .A(n319), .ZN(n309) );
  INV_X1 U226 ( .A(n318), .ZN(n306) );
  INV_X1 U227 ( .A(n318), .ZN(n308) );
  INV_X1 U228 ( .A(n318), .ZN(n307) );
  INV_X1 U229 ( .A(n320), .ZN(n314) );
  NAND2_X1 U230 ( .A1(n314), .A2(n377), .ZN(n380) );
  INV_X1 U231 ( .A(n319), .ZN(n312) );
  INV_X1 U232 ( .A(n319), .ZN(n313) );
  AND2_X1 U233 ( .A1(n257), .A2(n367), .ZN(n266) );
  INV_X1 U234 ( .A(n95), .ZN(n267) );
  NAND2_X1 U235 ( .A1(n348), .A2(n346), .ZN(n372) );
  NOR2_X1 U236 ( .A1(n372), .A2(n220), .ZN(n373) );
  CLKBUF_X1 U237 ( .A(n321), .Z(n320) );
  BUF_X1 U238 ( .A(n323), .Z(n316) );
  CLKBUF_X1 U239 ( .A(n322), .Z(n317) );
  CLKBUF_X1 U240 ( .A(n323), .Z(n315) );
  INV_X1 U241 ( .A(n160), .ZN(n341) );
  INV_X1 U242 ( .A(n129), .ZN(n321) );
  INV_X1 U243 ( .A(n129), .ZN(n322) );
  INV_X1 U244 ( .A(n129), .ZN(n323) );
  INV_X1 U245 ( .A(n90), .ZN(n327) );
  CLKBUF_X1 U246 ( .A(n62), .Z(n275) );
  XNOR2_X1 U247 ( .A(n370), .B(n344), .ZN(n62) );
  INV_X1 U248 ( .A(n273), .ZN(n324) );
  INV_X2 U249 ( .A(n217), .ZN(n326) );
  CLKBUF_X1 U250 ( .A(n280), .Z(n276) );
  NAND2_X1 U251 ( .A1(n380), .A2(n379), .ZN(n56) );
  XOR2_X1 U252 ( .A(n45), .B(n274), .Z(n352) );
  INV_X1 U253 ( .A(n64), .ZN(n277) );
  INV_X1 U254 ( .A(n277), .ZN(n278) );
  OR2_X1 U255 ( .A1(n374), .A2(n349), .ZN(n284) );
  CLKBUF_X1 U256 ( .A(n226), .Z(n281) );
  AND2_X2 U257 ( .A1(n376), .A2(n375), .ZN(n279) );
  AND2_X2 U258 ( .A1(n371), .A2(n232), .ZN(n280) );
  XNOR2_X1 U259 ( .A(n360), .B(n43), .ZN(n64) );
  OAI21_X1 U260 ( .B1(n240), .B2(n329), .A(n70), .ZN(n356) );
  INV_X1 U261 ( .A(n158), .ZN(n339) );
  NAND2_X1 U262 ( .A1(n374), .A2(n349), .ZN(n283) );
  NAND2_X2 U263 ( .A1(n283), .A2(n284), .ZN(n78) );
  OAI21_X1 U264 ( .B1(n370), .B2(n342), .A(n168), .ZN(n371) );
  INV_X1 U265 ( .A(n45), .ZN(n328) );
  NAND2_X1 U266 ( .A1(n369), .A2(n282), .ZN(n370) );
  INV_X1 U267 ( .A(n95), .ZN(n338) );
  INV_X1 U268 ( .A(n70), .ZN(n333) );
  NAND2_X1 U269 ( .A1(n354), .A2(n353), .ZN(n357) );
  INV_X1 U270 ( .A(n352), .ZN(n61) );
  NOR2_X1 U271 ( .A1(n364), .A2(n301), .ZN(n360) );
  NAND2_X1 U272 ( .A1(n300), .A2(n304), .ZN(n365) );
  NOR2_X1 U273 ( .A1(n365), .A2(n271), .ZN(n366) );
  NAND2_X1 U274 ( .A1(n328), .A2(n273), .ZN(n355) );
  OAI21_X1 U275 ( .B1(n232), .B2(n220), .A(n174), .ZN(n375) );
  NOR2_X1 U276 ( .A1(n365), .A2(n368), .ZN(n363) );
  INV_X2 U277 ( .A(n211), .ZN(n329) );
  INV_X2 U278 ( .A(n341), .ZN(n340) );
  INV_X2 U279 ( .A(n344), .ZN(n342) );
  INV_X1 U280 ( .A(n234), .ZN(n302) );
  INV_X1 U281 ( .A(n86), .ZN(n303) );
  INV_X1 U282 ( .A(n86), .ZN(n304) );
  INV_X1 U283 ( .A(n301), .ZN(n305) );
  INV_X1 U284 ( .A(n274), .ZN(n325) );
  INV_X1 U285 ( .A(n331), .ZN(n330) );
  INV_X1 U286 ( .A(n146), .ZN(n331) );
  INV_X1 U287 ( .A(n146), .ZN(n332) );
  INV_X1 U288 ( .A(n346), .ZN(n343) );
  INV_X1 U289 ( .A(n163), .ZN(n344) );
  INV_X1 U290 ( .A(n163), .ZN(n345) );
  INV_X1 U291 ( .A(n163), .ZN(n346) );
  INV_X1 U292 ( .A(n168), .ZN(n347) );
  INV_X1 U293 ( .A(n168), .ZN(n348) );
  INV_X1 U294 ( .A(n174), .ZN(n350) );
  INV_X1 U295 ( .A(n174), .ZN(n351) );
  INV_X1 U296 ( .A(n355), .ZN(n354) );
  NOR2_X1 U297 ( .A1(n330), .A2(n70), .ZN(n353) );
  NOR2_X1 U298 ( .A1(n330), .A2(n70), .ZN(n358) );
  NOR2_X1 U299 ( .A1(n70), .A2(n94), .ZN(n359) );
  NAND3_X1 U300 ( .A1(n268), .A2(n265), .A3(n359), .ZN(n364) );
  NOR2_X1 U301 ( .A1(n70), .A2(n94), .ZN(n362) );
  NOR2_X1 U302 ( .A1(n324), .A2(n45), .ZN(n361) );
  NAND3_X1 U303 ( .A1(n362), .A2(n361), .A3(n268), .ZN(n368) );
  NOR4_X1 U304 ( .A1(n231), .A2(n271), .A3(n43), .A4(n302), .ZN(n367) );
  NAND3_X1 U305 ( .A1(n254), .A2(n351), .A3(n373), .ZN(n376) );
  NAND2_X1 U306 ( .A1(n320), .A2(n376), .ZN(n379) );
  INV_X1 U307 ( .A(n379), .ZN(n381) );
  INV_X1 U308 ( .A(n376), .ZN(n377) );
  INV_X1 U309 ( .A(n380), .ZN(n378) );
endmodule


module Comparator_Nbit32 ( Diff, Cout, Sign, a, b, Ne, Eq, Gt, Ge, Lt, Le );
  input [31:0] Diff;
  input Cout, Sign, a, b;
  output Ne, Eq, Gt, Ge, Lt, Le;
  wire   n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;

  OR2_X1 U1 ( .A1(Diff[0]), .A2(Diff[1]), .ZN(n60) );
  NAND2_X1 U2 ( .A1(Ne), .A2(Ge), .ZN(Le) );
  NOR2_X1 U3 ( .A1(Diff[7]), .A2(Diff[6]), .ZN(n63) );
  XNOR2_X1 U4 ( .A(Cout), .B(n47), .ZN(Lt) );
  XNOR2_X1 U5 ( .A(a), .B(b), .ZN(n46) );
  INV_X1 U6 ( .A(Sign), .ZN(n45) );
  NOR2_X1 U7 ( .A1(n46), .A2(n45), .ZN(n47) );
  NOR2_X1 U8 ( .A1(Diff[27]), .A2(Diff[26]), .ZN(n49) );
  NOR2_X1 U9 ( .A1(Diff[25]), .A2(Diff[24]), .ZN(n48) );
  NAND2_X1 U10 ( .A1(n49), .A2(n48), .ZN(n53) );
  NOR2_X1 U11 ( .A1(Diff[31]), .A2(Diff[30]), .ZN(n51) );
  NOR2_X1 U12 ( .A1(Diff[29]), .A2(Diff[28]), .ZN(n50) );
  NAND2_X1 U13 ( .A1(n51), .A2(n50), .ZN(n52) );
  NOR2_X1 U14 ( .A1(n53), .A2(n52), .ZN(n71) );
  NOR2_X1 U15 ( .A1(Diff[19]), .A2(Diff[18]), .ZN(n55) );
  NOR2_X1 U16 ( .A1(Diff[17]), .A2(Diff[16]), .ZN(n54) );
  NAND2_X1 U17 ( .A1(n55), .A2(n54), .ZN(n59) );
  NOR2_X1 U18 ( .A1(Diff[23]), .A2(Diff[22]), .ZN(n57) );
  NOR2_X1 U19 ( .A1(Diff[21]), .A2(Diff[20]), .ZN(n56) );
  NAND2_X1 U20 ( .A1(n57), .A2(n56), .ZN(n58) );
  NOR2_X1 U21 ( .A1(n59), .A2(n58), .ZN(n70) );
  NOR2_X1 U22 ( .A1(Diff[5]), .A2(Diff[4]), .ZN(n62) );
  NOR3_X1 U23 ( .A1(n60), .A2(Diff[3]), .A3(Diff[2]), .ZN(n61) );
  NAND3_X1 U24 ( .A1(n63), .A2(n62), .A3(n61), .ZN(n68) );
  NOR2_X1 U25 ( .A1(Diff[15]), .A2(Diff[14]), .ZN(n66) );
  NOR2_X1 U26 ( .A1(Diff[13]), .A2(Diff[12]), .ZN(n65) );
  NOR4_X1 U27 ( .A1(Diff[9]), .A2(Diff[8]), .A3(Diff[11]), .A4(Diff[10]), .ZN(
        n64) );
  NAND3_X1 U28 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n67) );
  NOR2_X1 U29 ( .A1(n68), .A2(n67), .ZN(n69) );
  NAND3_X1 U30 ( .A1(n71), .A2(n70), .A3(n69), .ZN(Ne) );
  INV_X1 U31 ( .A(Lt), .ZN(Ge) );
  INV_X1 U32 ( .A(Le), .ZN(Gt) );
  INV_X1 U33 ( .A(Ne), .ZN(Eq) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE, 
        OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, n116, n117, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551;
  assign n116 = B[3];
  assign n117 = B[4];

  SHIFTER_GENERIC_N32_DW01_ash_0 C88 ( .A(A), .DATA_TC(1'b0), .SH({n117, n371, 
        B[2:0]}), .SH_TC(1'b0), .B({N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234}) );
  SHIFTER_GENERIC_N32_DW_sla_0 C86 ( .A(A), .SH({n117, n371, B[2:0]}), .SH_TC(
        1'b0), .B({N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202}) );
  SHIFTER_GENERIC_N32_DW_rash_0 C50 ( .A(A), .DATA_TC(1'b0), .SH({n117, n371, 
        B[2:0]}), .SH_TC(1'b0), .B({N168, N167, N166, N165, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137}) );
  SHIFTER_GENERIC_N32_DW_sra_0 C48 ( .A(A), .SH({n117, n371, B[2:0]}), .SH_TC(
        1'b0), .B({N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105}) );
  SHIFTER_GENERIC_N32_DW_lbsh_0 C10 ( .A(A), .SH({n117, n371, B[2:0]}), 
        .SH_TC(1'b0), .B({N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39}) );
  SHIFTER_GENERIC_N32_DW_rbsh_0 C8 ( .A(A), .SH({n117, n371, B[2:0]}), .SH_TC(
        1'b0), .B({N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7}) );
  AND2_X1 U1 ( .A1(N240), .A2(n368), .ZN(n323) );
  AND2_X1 U2 ( .A1(N241), .A2(n368), .ZN(n324) );
  AND2_X1 U3 ( .A1(N239), .A2(n368), .ZN(n325) );
  AND2_X1 U4 ( .A1(N238), .A2(n368), .ZN(n326) );
  AND2_X1 U5 ( .A1(N151), .A2(n359), .ZN(n327) );
  AND2_X1 U6 ( .A1(N160), .A2(n358), .ZN(n328) );
  AND2_X1 U7 ( .A1(N105), .A2(n360), .ZN(n329) );
  AND2_X1 U8 ( .A1(N106), .A2(n360), .ZN(n330) );
  AND2_X1 U9 ( .A1(N107), .A2(n360), .ZN(n331) );
  AND2_X1 U10 ( .A1(N116), .A2(n360), .ZN(n332) );
  AND2_X1 U11 ( .A1(N117), .A2(n360), .ZN(n333) );
  AND2_X1 U12 ( .A1(N121), .A2(n361), .ZN(n334) );
  AND2_X1 U13 ( .A1(N147), .A2(n358), .ZN(n335) );
  AND2_X1 U14 ( .A1(N150), .A2(n359), .ZN(n336) );
  AND2_X1 U15 ( .A1(N152), .A2(n359), .ZN(n337) );
  AND2_X1 U16 ( .A1(N156), .A2(n359), .ZN(n338) );
  AND2_X1 U17 ( .A1(N157), .A2(n359), .ZN(n339) );
  AND2_X1 U18 ( .A1(N158), .A2(n359), .ZN(n340) );
  AND2_X1 U19 ( .A1(N159), .A2(n359), .ZN(n341) );
  AND2_X1 U20 ( .A1(N119), .A2(n361), .ZN(n342) );
  AND2_X1 U21 ( .A1(N128), .A2(n361), .ZN(n343) );
  AND2_X1 U22 ( .A1(N129), .A2(n361), .ZN(n344) );
  CLKBUF_X1 U23 ( .A(n116), .Z(n371) );
  BUF_X1 U24 ( .A(n347), .Z(n370) );
  BUF_X1 U25 ( .A(n348), .Z(n366) );
  BUF_X1 U26 ( .A(n347), .Z(n369) );
  BUF_X1 U27 ( .A(n348), .Z(n365) );
  BUF_X1 U28 ( .A(n508), .Z(n360) );
  BUF_X1 U29 ( .A(n508), .Z(n361) );
  AND2_X1 U30 ( .A1(n480), .A2(n345), .ZN(n483) );
  AND2_X1 U31 ( .A1(n482), .A2(n481), .ZN(n345) );
  AND2_X1 U32 ( .A1(n473), .A2(n346), .ZN(n476) );
  AND2_X1 U33 ( .A1(n475), .A2(n474), .ZN(n346) );
  BUF_X1 U34 ( .A(n357), .Z(n363) );
  BUF_X1 U35 ( .A(n547), .Z(n367) );
  BUF_X1 U36 ( .A(n357), .Z(n364) );
  BUF_X1 U37 ( .A(n547), .Z(n368) );
  BUF_X1 U38 ( .A(n503), .Z(n358) );
  BUF_X1 U39 ( .A(n503), .Z(n359) );
  NAND4_X1 U40 ( .A1(n531), .A2(n530), .A3(n529), .A4(n528), .ZN(OUTPUT[27])
         );
  NAND2_X1 U41 ( .A1(N66), .A2(n365), .ZN(n529) );
  AOI22_X1 U42 ( .A1(N132), .A2(n527), .B1(N164), .B2(n546), .ZN(n531) );
  AOI22_X1 U43 ( .A1(N34), .A2(n369), .B1(N261), .B2(n367), .ZN(n528) );
  NAND4_X1 U44 ( .A1(n551), .A2(n550), .A3(n549), .A4(n548), .ZN(OUTPUT[31])
         );
  NAND2_X1 U45 ( .A1(N70), .A2(n365), .ZN(n549) );
  AOI22_X1 U46 ( .A1(N136), .A2(n527), .B1(N168), .B2(n546), .ZN(n551) );
  AOI22_X1 U47 ( .A1(N38), .A2(n369), .B1(N265), .B2(n367), .ZN(n548) );
  NAND4_X1 U48 ( .A1(n535), .A2(n534), .A3(n533), .A4(n532), .ZN(OUTPUT[28])
         );
  NAND2_X1 U49 ( .A1(N67), .A2(n365), .ZN(n533) );
  AOI22_X1 U50 ( .A1(N133), .A2(n527), .B1(N165), .B2(n546), .ZN(n535) );
  AOI22_X1 U51 ( .A1(N35), .A2(n369), .B1(N262), .B2(n367), .ZN(n532) );
  NAND4_X1 U52 ( .A1(n543), .A2(n542), .A3(n541), .A4(n540), .ZN(OUTPUT[30])
         );
  NAND2_X1 U53 ( .A1(N69), .A2(n365), .ZN(n541) );
  AOI22_X1 U54 ( .A1(N135), .A2(n527), .B1(N167), .B2(n546), .ZN(n543) );
  AOI22_X1 U55 ( .A1(N37), .A2(n369), .B1(N264), .B2(n367), .ZN(n540) );
  NAND4_X1 U56 ( .A1(n526), .A2(n525), .A3(n524), .A4(n523), .ZN(OUTPUT[26])
         );
  NAND2_X1 U57 ( .A1(N65), .A2(n365), .ZN(n524) );
  AOI22_X1 U58 ( .A1(N131), .A2(n527), .B1(N163), .B2(n546), .ZN(n526) );
  AOI22_X1 U59 ( .A1(N33), .A2(n369), .B1(N260), .B2(n367), .ZN(n523) );
  NAND4_X1 U60 ( .A1(n539), .A2(n538), .A3(n537), .A4(n536), .ZN(OUTPUT[29])
         );
  NAND2_X1 U61 ( .A1(N68), .A2(n365), .ZN(n537) );
  AOI22_X1 U62 ( .A1(N134), .A2(n527), .B1(N166), .B2(n546), .ZN(n539) );
  AOI22_X1 U63 ( .A1(N36), .A2(n369), .B1(N263), .B2(n367), .ZN(n536) );
  INV_X1 U64 ( .A(n544), .ZN(n527) );
  AND2_X1 U65 ( .A1(n374), .A2(n376), .ZN(n347) );
  AND2_X1 U66 ( .A1(n374), .A2(LEFT_RIGHT), .ZN(n348) );
  NAND2_X1 U67 ( .A1(N229), .A2(n363), .ZN(n530) );
  NAND2_X1 U68 ( .A1(N228), .A2(n363), .ZN(n525) );
  NAND2_X1 U69 ( .A1(N233), .A2(n363), .ZN(n550) );
  NAND2_X1 U70 ( .A1(N230), .A2(n363), .ZN(n534) );
  NAND2_X1 U71 ( .A1(N232), .A2(n363), .ZN(n542) );
  NAND2_X1 U72 ( .A1(N231), .A2(n363), .ZN(n538) );
  AND2_X1 U73 ( .A1(N243), .A2(n368), .ZN(n349) );
  AND2_X1 U74 ( .A1(N244), .A2(n368), .ZN(n350) );
  AND2_X1 U75 ( .A1(N242), .A2(n368), .ZN(n351) );
  AND2_X1 U76 ( .A1(N245), .A2(n368), .ZN(n352) );
  AND2_X1 U77 ( .A1(N247), .A2(n368), .ZN(n353) );
  AND2_X1 U78 ( .A1(N249), .A2(n368), .ZN(n354) );
  AND2_X1 U79 ( .A1(N248), .A2(n368), .ZN(n355) );
  AND2_X1 U80 ( .A1(N246), .A2(n368), .ZN(n356) );
  NOR2_X1 U81 ( .A1(n545), .A2(n516), .ZN(n517) );
  NOR2_X1 U82 ( .A1(n408), .A2(n384), .ZN(n385) );
  NOR2_X1 U83 ( .A1(n408), .A2(n372), .ZN(n373) );
  INV_X1 U84 ( .A(n545), .ZN(n546) );
  AND3_X1 U85 ( .A1(SHIFT_ROTATE), .A2(LEFT_RIGHT), .A3(n377), .ZN(n357) );
  NAND3_X1 U86 ( .A1(LOGIC_ARITH), .A2(SHIFT_ROTATE), .A3(n376), .ZN(n545) );
  CLKBUF_X1 U87 ( .A(n508), .Z(n362) );
  INV_X1 U88 ( .A(SHIFT_ROTATE), .ZN(n374) );
  INV_X1 U89 ( .A(LEFT_RIGHT), .ZN(n376) );
  NAND3_X1 U90 ( .A1(LOGIC_ARITH), .A2(LEFT_RIGHT), .A3(SHIFT_ROTATE), .ZN(
        n408) );
  INV_X1 U91 ( .A(N234), .ZN(n372) );
  AOI21_X1 U92 ( .B1(N7), .B2(n369), .A(n373), .ZN(n383) );
  NAND2_X1 U93 ( .A1(N39), .A2(n366), .ZN(n382) );
  INV_X1 U94 ( .A(LOGIC_ARITH), .ZN(n377) );
  NOR2_X1 U95 ( .A1(LEFT_RIGHT), .A2(n374), .ZN(n375) );
  NAND2_X1 U96 ( .A1(n377), .A2(n375), .ZN(n544) );
  INV_X1 U97 ( .A(n544), .ZN(n508) );
  INV_X1 U98 ( .A(n545), .ZN(n503) );
  NAND2_X1 U99 ( .A1(N137), .A2(n358), .ZN(n379) );
  NAND2_X1 U100 ( .A1(N202), .A2(n364), .ZN(n378) );
  NAND2_X1 U101 ( .A1(n379), .A2(n378), .ZN(n380) );
  NOR2_X1 U102 ( .A1(n329), .A2(n380), .ZN(n381) );
  NAND3_X1 U103 ( .A1(n383), .A2(n382), .A3(n381), .ZN(OUTPUT[0]) );
  INV_X1 U104 ( .A(N235), .ZN(n384) );
  AOI21_X1 U105 ( .B1(N8), .B2(n369), .A(n385), .ZN(n391) );
  NAND2_X1 U106 ( .A1(N40), .A2(n366), .ZN(n390) );
  NAND2_X1 U107 ( .A1(N138), .A2(n358), .ZN(n387) );
  NAND2_X1 U108 ( .A1(N203), .A2(n364), .ZN(n386) );
  NAND2_X1 U109 ( .A1(n387), .A2(n386), .ZN(n388) );
  NOR2_X1 U110 ( .A1(n330), .A2(n388), .ZN(n389) );
  NAND3_X1 U111 ( .A1(n391), .A2(n390), .A3(n389), .ZN(OUTPUT[1]) );
  INV_X1 U112 ( .A(N236), .ZN(n392) );
  NOR2_X1 U113 ( .A1(n408), .A2(n392), .ZN(n393) );
  AOI21_X1 U114 ( .B1(N9), .B2(n370), .A(n393), .ZN(n399) );
  NAND2_X1 U115 ( .A1(N41), .A2(n366), .ZN(n398) );
  NAND2_X1 U116 ( .A1(N139), .A2(n358), .ZN(n395) );
  NAND2_X1 U117 ( .A1(N204), .A2(n364), .ZN(n394) );
  NAND2_X1 U118 ( .A1(n395), .A2(n394), .ZN(n396) );
  NOR2_X1 U119 ( .A1(n331), .A2(n396), .ZN(n397) );
  NAND3_X1 U120 ( .A1(n399), .A2(n398), .A3(n397), .ZN(OUTPUT[2]) );
  INV_X1 U121 ( .A(N237), .ZN(n400) );
  NOR2_X1 U122 ( .A1(n408), .A2(n400), .ZN(n401) );
  AOI21_X1 U123 ( .B1(N10), .B2(n370), .A(n401), .ZN(n407) );
  NAND2_X1 U124 ( .A1(N42), .A2(n366), .ZN(n406) );
  NAND2_X1 U125 ( .A1(N140), .A2(n358), .ZN(n403) );
  NAND2_X1 U126 ( .A1(N205), .A2(n364), .ZN(n402) );
  NAND2_X1 U127 ( .A1(n403), .A2(n402), .ZN(n404) );
  AOI21_X1 U128 ( .B1(N108), .B2(n360), .A(n404), .ZN(n405) );
  NAND3_X1 U129 ( .A1(n407), .A2(n406), .A3(n405), .ZN(OUTPUT[3]) );
  INV_X1 U130 ( .A(n408), .ZN(n547) );
  AOI21_X1 U131 ( .B1(N11), .B2(n370), .A(n326), .ZN(n414) );
  NAND2_X1 U132 ( .A1(N43), .A2(n366), .ZN(n413) );
  NAND2_X1 U133 ( .A1(N141), .A2(n358), .ZN(n410) );
  NAND2_X1 U134 ( .A1(N206), .A2(n364), .ZN(n409) );
  NAND2_X1 U135 ( .A1(n410), .A2(n409), .ZN(n411) );
  AOI21_X1 U136 ( .B1(N109), .B2(n360), .A(n411), .ZN(n412) );
  NAND3_X1 U137 ( .A1(n414), .A2(n413), .A3(n412), .ZN(OUTPUT[4]) );
  AOI21_X1 U138 ( .B1(N12), .B2(n370), .A(n325), .ZN(n420) );
  NAND2_X1 U139 ( .A1(N44), .A2(n366), .ZN(n419) );
  NAND2_X1 U140 ( .A1(N142), .A2(n358), .ZN(n416) );
  NAND2_X1 U141 ( .A1(N207), .A2(n364), .ZN(n415) );
  NAND2_X1 U142 ( .A1(n416), .A2(n415), .ZN(n417) );
  AOI21_X1 U143 ( .B1(N110), .B2(n360), .A(n417), .ZN(n418) );
  NAND3_X1 U144 ( .A1(n420), .A2(n419), .A3(n418), .ZN(OUTPUT[5]) );
  AOI21_X1 U145 ( .B1(N13), .B2(n370), .A(n323), .ZN(n426) );
  NAND2_X1 U146 ( .A1(N45), .A2(n366), .ZN(n425) );
  NAND2_X1 U147 ( .A1(N143), .A2(n358), .ZN(n422) );
  NAND2_X1 U148 ( .A1(N208), .A2(n364), .ZN(n421) );
  NAND2_X1 U149 ( .A1(n422), .A2(n421), .ZN(n423) );
  AOI21_X1 U150 ( .B1(N111), .B2(n360), .A(n423), .ZN(n424) );
  NAND3_X1 U151 ( .A1(n426), .A2(n425), .A3(n424), .ZN(OUTPUT[6]) );
  AOI21_X1 U152 ( .B1(N14), .B2(n370), .A(n324), .ZN(n432) );
  NAND2_X1 U153 ( .A1(N46), .A2(n366), .ZN(n431) );
  NAND2_X1 U154 ( .A1(N144), .A2(n358), .ZN(n428) );
  NAND2_X1 U155 ( .A1(N209), .A2(n364), .ZN(n427) );
  NAND2_X1 U156 ( .A1(n428), .A2(n427), .ZN(n429) );
  AOI21_X1 U157 ( .B1(N112), .B2(n360), .A(n429), .ZN(n430) );
  NAND3_X1 U158 ( .A1(n432), .A2(n431), .A3(n430), .ZN(OUTPUT[7]) );
  AOI21_X1 U159 ( .B1(N15), .B2(n369), .A(n351), .ZN(n438) );
  NAND2_X1 U160 ( .A1(N47), .A2(n366), .ZN(n437) );
  NAND2_X1 U161 ( .A1(N145), .A2(n358), .ZN(n434) );
  NAND2_X1 U162 ( .A1(N210), .A2(n364), .ZN(n433) );
  NAND2_X1 U163 ( .A1(n434), .A2(n433), .ZN(n435) );
  AOI21_X1 U164 ( .B1(N113), .B2(n360), .A(n435), .ZN(n436) );
  NAND3_X1 U165 ( .A1(n438), .A2(n437), .A3(n436), .ZN(OUTPUT[8]) );
  AOI21_X1 U166 ( .B1(N16), .B2(n369), .A(n349), .ZN(n441) );
  NAND2_X1 U167 ( .A1(N48), .A2(n366), .ZN(n440) );
  AOI222_X1 U168 ( .A1(N114), .A2(n360), .B1(N211), .B2(n364), .C1(N146), .C2(
        n359), .ZN(n439) );
  NAND3_X1 U169 ( .A1(n441), .A2(n440), .A3(n439), .ZN(OUTPUT[9]) );
  AOI21_X1 U170 ( .B1(N17), .B2(n369), .A(n350), .ZN(n444) );
  NAND2_X1 U171 ( .A1(N49), .A2(n366), .ZN(n443) );
  AOI221_X1 U172 ( .B1(N115), .B2(n362), .C1(N212), .C2(n363), .A(n335), .ZN(
        n442) );
  NAND3_X1 U173 ( .A1(n444), .A2(n443), .A3(n442), .ZN(OUTPUT[10]) );
  AOI21_X1 U174 ( .B1(N18), .B2(n369), .A(n352), .ZN(n450) );
  NAND2_X1 U175 ( .A1(N50), .A2(n366), .ZN(n449) );
  NAND2_X1 U176 ( .A1(N148), .A2(n358), .ZN(n446) );
  NAND2_X1 U177 ( .A1(N213), .A2(n364), .ZN(n445) );
  NAND2_X1 U178 ( .A1(n446), .A2(n445), .ZN(n447) );
  NOR2_X1 U179 ( .A1(n332), .A2(n447), .ZN(n448) );
  NAND3_X1 U180 ( .A1(n450), .A2(n449), .A3(n448), .ZN(OUTPUT[11]) );
  AOI21_X1 U181 ( .B1(N19), .B2(n369), .A(n356), .ZN(n456) );
  NAND2_X1 U182 ( .A1(N51), .A2(n366), .ZN(n455) );
  NAND2_X1 U183 ( .A1(N149), .A2(n359), .ZN(n452) );
  NAND2_X1 U184 ( .A1(N214), .A2(n364), .ZN(n451) );
  NAND2_X1 U185 ( .A1(n452), .A2(n451), .ZN(n453) );
  NOR2_X1 U186 ( .A1(n333), .A2(n453), .ZN(n454) );
  NAND3_X1 U187 ( .A1(n456), .A2(n455), .A3(n454), .ZN(OUTPUT[12]) );
  AOI21_X1 U188 ( .B1(N20), .B2(n369), .A(n353), .ZN(n459) );
  NAND2_X1 U189 ( .A1(N52), .A2(n366), .ZN(n458) );
  AOI221_X1 U190 ( .B1(N118), .B2(n361), .C1(N215), .C2(n363), .A(n336), .ZN(
        n457) );
  NAND3_X1 U191 ( .A1(n459), .A2(n458), .A3(n457), .ZN(OUTPUT[13]) );
  AOI21_X1 U192 ( .B1(N21), .B2(n369), .A(n355), .ZN(n462) );
  NAND2_X1 U193 ( .A1(N53), .A2(n366), .ZN(n461) );
  AOI211_X1 U194 ( .C1(N216), .C2(n364), .A(n342), .B(n327), .ZN(n460) );
  NAND3_X1 U195 ( .A1(n462), .A2(n461), .A3(n460), .ZN(OUTPUT[14]) );
  AOI21_X1 U196 ( .B1(N22), .B2(n369), .A(n354), .ZN(n465) );
  NAND2_X1 U197 ( .A1(N54), .A2(n366), .ZN(n464) );
  AOI221_X1 U198 ( .B1(N120), .B2(n361), .C1(N217), .C2(n363), .A(n337), .ZN(
        n463) );
  NAND3_X1 U199 ( .A1(n465), .A2(n464), .A3(n463), .ZN(OUTPUT[15]) );
  NAND2_X1 U200 ( .A1(N23), .A2(n370), .ZN(n472) );
  NAND2_X1 U201 ( .A1(N250), .A2(n367), .ZN(n471) );
  NAND2_X1 U202 ( .A1(N55), .A2(n365), .ZN(n470) );
  NAND2_X1 U203 ( .A1(N153), .A2(n359), .ZN(n467) );
  NAND2_X1 U204 ( .A1(N218), .A2(n364), .ZN(n466) );
  NAND2_X1 U205 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U206 ( .A1(n334), .A2(n468), .ZN(n469) );
  NAND4_X1 U207 ( .A1(n472), .A2(n471), .A3(n470), .A4(n469), .ZN(OUTPUT[16])
         );
  NAND2_X1 U208 ( .A1(N24), .A2(n370), .ZN(n479) );
  NAND2_X1 U209 ( .A1(N251), .A2(n367), .ZN(n478) );
  NAND2_X1 U210 ( .A1(N56), .A2(n365), .ZN(n477) );
  NAND2_X1 U211 ( .A1(N122), .A2(n361), .ZN(n473) );
  NAND2_X1 U212 ( .A1(N154), .A2(n359), .ZN(n475) );
  NAND2_X1 U213 ( .A1(N219), .A2(n364), .ZN(n474) );
  NAND4_X1 U214 ( .A1(n479), .A2(n478), .A3(n477), .A4(n476), .ZN(OUTPUT[17])
         );
  NAND2_X1 U215 ( .A1(N25), .A2(n370), .ZN(n486) );
  NAND2_X1 U216 ( .A1(N252), .A2(n367), .ZN(n485) );
  NAND2_X1 U217 ( .A1(N57), .A2(n365), .ZN(n484) );
  NAND2_X1 U218 ( .A1(N123), .A2(n361), .ZN(n480) );
  NAND2_X1 U219 ( .A1(N155), .A2(n359), .ZN(n482) );
  NAND2_X1 U220 ( .A1(N220), .A2(n364), .ZN(n481) );
  NAND4_X1 U221 ( .A1(n486), .A2(n485), .A3(n484), .A4(n483), .ZN(OUTPUT[18])
         );
  NAND2_X1 U222 ( .A1(N26), .A2(n370), .ZN(n490) );
  NAND2_X1 U223 ( .A1(N253), .A2(n367), .ZN(n489) );
  NAND2_X1 U224 ( .A1(N58), .A2(n365), .ZN(n488) );
  AOI221_X1 U225 ( .B1(N124), .B2(n361), .C1(N221), .C2(n363), .A(n338), .ZN(
        n487) );
  NAND4_X1 U226 ( .A1(n490), .A2(n489), .A3(n488), .A4(n487), .ZN(OUTPUT[19])
         );
  NAND2_X1 U227 ( .A1(N27), .A2(n370), .ZN(n494) );
  NAND2_X1 U228 ( .A1(N254), .A2(n367), .ZN(n493) );
  NAND2_X1 U229 ( .A1(N59), .A2(n365), .ZN(n492) );
  AOI221_X1 U230 ( .B1(N125), .B2(n361), .C1(N222), .C2(n363), .A(n339), .ZN(
        n491) );
  NAND4_X1 U231 ( .A1(n494), .A2(n493), .A3(n492), .A4(n491), .ZN(OUTPUT[20])
         );
  NAND2_X1 U232 ( .A1(N28), .A2(n370), .ZN(n498) );
  NAND2_X1 U233 ( .A1(N255), .A2(n367), .ZN(n497) );
  NAND2_X1 U234 ( .A1(N60), .A2(n365), .ZN(n496) );
  AOI221_X1 U235 ( .B1(N126), .B2(n361), .C1(N223), .C2(n363), .A(n340), .ZN(
        n495) );
  NAND4_X1 U236 ( .A1(n498), .A2(n497), .A3(n496), .A4(n495), .ZN(OUTPUT[21])
         );
  NAND2_X1 U237 ( .A1(N29), .A2(n370), .ZN(n502) );
  NAND2_X1 U238 ( .A1(N256), .A2(n367), .ZN(n501) );
  NAND2_X1 U239 ( .A1(N61), .A2(n365), .ZN(n500) );
  AOI221_X1 U240 ( .B1(N127), .B2(n361), .C1(N224), .C2(n363), .A(n341), .ZN(
        n499) );
  NAND4_X1 U241 ( .A1(n502), .A2(n501), .A3(n500), .A4(n499), .ZN(OUTPUT[22])
         );
  NAND2_X1 U242 ( .A1(N30), .A2(n370), .ZN(n507) );
  NAND2_X1 U243 ( .A1(N257), .A2(n367), .ZN(n506) );
  NAND2_X1 U244 ( .A1(N62), .A2(n365), .ZN(n505) );
  AOI211_X1 U245 ( .C1(N225), .C2(n363), .A(n343), .B(n328), .ZN(n504) );
  NAND4_X1 U246 ( .A1(n507), .A2(n506), .A3(n505), .A4(n504), .ZN(OUTPUT[23])
         );
  NAND2_X1 U247 ( .A1(N31), .A2(n370), .ZN(n514) );
  NAND2_X1 U248 ( .A1(N258), .A2(n367), .ZN(n513) );
  NAND2_X1 U249 ( .A1(N63), .A2(n365), .ZN(n512) );
  INV_X1 U250 ( .A(N161), .ZN(n509) );
  NOR2_X1 U251 ( .A1(n545), .A2(n509), .ZN(n510) );
  AOI211_X1 U252 ( .C1(N226), .C2(n363), .A(n344), .B(n510), .ZN(n511) );
  NAND4_X1 U253 ( .A1(n514), .A2(n513), .A3(n512), .A4(n511), .ZN(OUTPUT[24])
         );
  NAND2_X1 U254 ( .A1(N32), .A2(n370), .ZN(n522) );
  NAND2_X1 U255 ( .A1(N259), .A2(n367), .ZN(n521) );
  NAND2_X1 U256 ( .A1(N64), .A2(n365), .ZN(n520) );
  INV_X1 U257 ( .A(N130), .ZN(n515) );
  NOR2_X1 U258 ( .A1(n544), .A2(n515), .ZN(n518) );
  INV_X1 U259 ( .A(N162), .ZN(n516) );
  AOI211_X1 U260 ( .C1(N227), .C2(n363), .A(n518), .B(n517), .ZN(n519) );
  NAND4_X1 U261 ( .A1(n522), .A2(n521), .A3(n520), .A4(n519), .ZN(OUTPUT[25])
         );
endmodule


module Add_gen_N32 ( A, B, sub, S, Co, Sign_OF, Unsign_OF );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input sub;
  output Co, Sign_OF, Unsign_OF;
  wire   n3, n8, n9, n10, n11, n12;
  wire   [31:0] BS;
  assign n3 = sub;

  xor_gen_N32_1 SUBTR ( .A(B), .B({n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, 
        n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, n8, 
        n8, n8, n8}), .C(BS) );
  p4adder_N32_0 ADDER ( .A(A), .B(BS), .Cin(n8), .S(S), .Cout(Co) );
  INV_X1 U1 ( .A(n3), .ZN(n9) );
  XNOR2_X1 U2 ( .A(n12), .B(n11), .ZN(Sign_OF) );
  INV_X4 U3 ( .A(n9), .ZN(n8) );
  XNOR2_X1 U4 ( .A(Co), .B(n9), .ZN(Unsign_OF) );
  INV_X1 U5 ( .A(BS[31]), .ZN(n10) );
  XNOR2_X1 U6 ( .A(S[31]), .B(n10), .ZN(n12) );
  XNOR2_X1 U7 ( .A(A[31]), .B(Co), .ZN(n11) );
endmodule


module xor_gen_N32_0 ( A, B, C );
  input [31:0] A;
  input [31:0] B;
  output [31:0] C;
  wire   n1, n2, n3;

  XNOR2_X1 U1 ( .A(A[2]), .B(n3), .ZN(C[2]) );
  XNOR2_X1 U2 ( .A(A[0]), .B(n1), .ZN(C[0]) );
  XNOR2_X1 U3 ( .A(A[1]), .B(n2), .ZN(C[1]) );
  INV_X1 U4 ( .A(B[0]), .ZN(n1) );
  INV_X1 U5 ( .A(B[1]), .ZN(n2) );
  INV_X1 U6 ( .A(B[2]), .ZN(n3) );
  XOR2_X1 U7 ( .A(A[3]), .B(B[3]), .Z(C[3]) );
  XOR2_X1 U8 ( .A(A[4]), .B(B[4]), .Z(C[4]) );
  XOR2_X1 U9 ( .A(A[5]), .B(B[5]), .Z(C[5]) );
  XOR2_X1 U10 ( .A(A[6]), .B(B[6]), .Z(C[6]) );
  XOR2_X1 U11 ( .A(A[7]), .B(B[7]), .Z(C[7]) );
  XOR2_X1 U12 ( .A(A[8]), .B(B[8]), .Z(C[8]) );
  XOR2_X1 U13 ( .A(A[9]), .B(B[9]), .Z(C[9]) );
  XOR2_X1 U14 ( .A(A[10]), .B(B[10]), .Z(C[10]) );
  XOR2_X1 U15 ( .A(A[11]), .B(B[11]), .Z(C[11]) );
  XOR2_X1 U16 ( .A(A[12]), .B(B[12]), .Z(C[12]) );
  XOR2_X1 U17 ( .A(A[13]), .B(B[13]), .Z(C[13]) );
  XOR2_X1 U18 ( .A(A[14]), .B(B[14]), .Z(C[14]) );
  XOR2_X1 U19 ( .A(A[15]), .B(B[15]), .Z(C[15]) );
  XOR2_X1 U20 ( .A(A[16]), .B(B[16]), .Z(C[16]) );
  XOR2_X1 U21 ( .A(A[17]), .B(B[17]), .Z(C[17]) );
  XOR2_X1 U22 ( .A(A[18]), .B(B[18]), .Z(C[18]) );
  XOR2_X1 U23 ( .A(A[19]), .B(B[19]), .Z(C[19]) );
  XOR2_X1 U24 ( .A(A[20]), .B(B[20]), .Z(C[20]) );
  XOR2_X1 U25 ( .A(A[21]), .B(B[21]), .Z(C[21]) );
  XOR2_X1 U26 ( .A(A[22]), .B(B[22]), .Z(C[22]) );
  XOR2_X1 U27 ( .A(A[23]), .B(B[23]), .Z(C[23]) );
  XOR2_X1 U28 ( .A(A[24]), .B(B[24]), .Z(C[24]) );
  XOR2_X1 U29 ( .A(A[25]), .B(B[25]), .Z(C[25]) );
  XOR2_X1 U30 ( .A(A[26]), .B(B[26]), .Z(C[26]) );
  XOR2_X1 U31 ( .A(A[27]), .B(B[27]), .Z(C[27]) );
  XOR2_X1 U32 ( .A(A[28]), .B(B[28]), .Z(C[28]) );
  XOR2_X1 U33 ( .A(A[29]), .B(B[29]), .Z(C[29]) );
  XOR2_X1 U34 ( .A(A[30]), .B(B[30]), .Z(C[30]) );
  XOR2_X1 U35 ( .A(A[31]), .B(B[31]), .Z(C[31]) );
endmodule


module or_gen_N32 ( A, B, C );
  input [31:0] A;
  input [31:0] B;
  output [31:0] C;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126;

  OR2_X1 U1 ( .A1(B[15]), .A2(A[15]), .ZN(C[15]) );
  INV_X1 U2 ( .A(A[7]), .ZN(n65) );
  INV_X1 U3 ( .A(A[6]), .ZN(n66) );
  INV_X1 U4 ( .A(B[0]), .ZN(n67) );
  INV_X1 U5 ( .A(B[1]), .ZN(n68) );
  INV_X1 U6 ( .A(B[2]), .ZN(n69) );
  INV_X1 U7 ( .A(B[3]), .ZN(n70) );
  INV_X1 U8 ( .A(A[0]), .ZN(n71) );
  INV_X1 U9 ( .A(A[1]), .ZN(n72) );
  INV_X1 U10 ( .A(A[2]), .ZN(n73) );
  INV_X1 U11 ( .A(A[3]), .ZN(n74) );
  INV_X1 U12 ( .A(A[4]), .ZN(n75) );
  INV_X1 U13 ( .A(A[5]), .ZN(n76) );
  INV_X1 U14 ( .A(A[8]), .ZN(n77) );
  INV_X1 U15 ( .A(A[9]), .ZN(n78) );
  INV_X1 U16 ( .A(A[10]), .ZN(n79) );
  INV_X1 U17 ( .A(A[11]), .ZN(n80) );
  INV_X1 U18 ( .A(A[12]), .ZN(n81) );
  INV_X1 U19 ( .A(A[13]), .ZN(n82) );
  INV_X1 U20 ( .A(A[14]), .ZN(n83) );
  INV_X1 U21 ( .A(A[20]), .ZN(n84) );
  INV_X1 U22 ( .A(A[22]), .ZN(n85) );
  INV_X1 U23 ( .A(A[24]), .ZN(n86) );
  INV_X1 U24 ( .A(A[25]), .ZN(n87) );
  INV_X1 U25 ( .A(A[26]), .ZN(n88) );
  NAND2_X1 U26 ( .A1(n67), .A2(n71), .ZN(C[0]) );
  NAND2_X1 U27 ( .A1(n68), .A2(n72), .ZN(C[1]) );
  NAND2_X1 U28 ( .A1(n69), .A2(n73), .ZN(C[2]) );
  NAND2_X1 U29 ( .A1(n70), .A2(n74), .ZN(C[3]) );
  INV_X1 U30 ( .A(B[4]), .ZN(n89) );
  NAND2_X1 U31 ( .A1(n89), .A2(n75), .ZN(C[4]) );
  INV_X1 U32 ( .A(B[5]), .ZN(n90) );
  NAND2_X1 U33 ( .A1(n90), .A2(n76), .ZN(C[5]) );
  INV_X1 U34 ( .A(B[6]), .ZN(n91) );
  NAND2_X1 U35 ( .A1(n91), .A2(n66), .ZN(C[6]) );
  INV_X1 U36 ( .A(B[7]), .ZN(n92) );
  NAND2_X1 U37 ( .A1(n92), .A2(n65), .ZN(C[7]) );
  INV_X1 U38 ( .A(B[8]), .ZN(n93) );
  NAND2_X1 U39 ( .A1(n93), .A2(n77), .ZN(C[8]) );
  INV_X1 U40 ( .A(B[9]), .ZN(n94) );
  NAND2_X1 U41 ( .A1(n94), .A2(n78), .ZN(C[9]) );
  INV_X1 U42 ( .A(B[10]), .ZN(n95) );
  NAND2_X1 U43 ( .A1(n95), .A2(n79), .ZN(C[10]) );
  INV_X1 U44 ( .A(B[11]), .ZN(n96) );
  NAND2_X1 U45 ( .A1(n96), .A2(n80), .ZN(C[11]) );
  INV_X1 U46 ( .A(B[12]), .ZN(n97) );
  NAND2_X1 U47 ( .A1(n97), .A2(n81), .ZN(C[12]) );
  INV_X1 U48 ( .A(B[13]), .ZN(n98) );
  NAND2_X1 U49 ( .A1(n98), .A2(n82), .ZN(C[13]) );
  INV_X1 U50 ( .A(B[14]), .ZN(n99) );
  NAND2_X1 U51 ( .A1(n99), .A2(n83), .ZN(C[14]) );
  INV_X1 U52 ( .A(B[16]), .ZN(n101) );
  INV_X1 U53 ( .A(A[16]), .ZN(n100) );
  NAND2_X1 U54 ( .A1(n101), .A2(n100), .ZN(C[16]) );
  INV_X1 U55 ( .A(B[17]), .ZN(n103) );
  INV_X1 U56 ( .A(A[17]), .ZN(n102) );
  NAND2_X1 U57 ( .A1(n103), .A2(n102), .ZN(C[17]) );
  INV_X1 U58 ( .A(B[18]), .ZN(n105) );
  INV_X1 U59 ( .A(A[18]), .ZN(n104) );
  NAND2_X1 U60 ( .A1(n105), .A2(n104), .ZN(C[18]) );
  INV_X1 U61 ( .A(B[19]), .ZN(n107) );
  INV_X1 U62 ( .A(A[19]), .ZN(n106) );
  NAND2_X1 U63 ( .A1(n107), .A2(n106), .ZN(C[19]) );
  INV_X1 U64 ( .A(B[20]), .ZN(n108) );
  NAND2_X1 U65 ( .A1(n108), .A2(n84), .ZN(C[20]) );
  INV_X1 U66 ( .A(B[21]), .ZN(n110) );
  INV_X1 U67 ( .A(A[21]), .ZN(n109) );
  NAND2_X1 U68 ( .A1(n110), .A2(n109), .ZN(C[21]) );
  INV_X1 U69 ( .A(B[22]), .ZN(n111) );
  NAND2_X1 U70 ( .A1(n111), .A2(n85), .ZN(C[22]) );
  INV_X1 U71 ( .A(B[23]), .ZN(n113) );
  INV_X1 U72 ( .A(A[23]), .ZN(n112) );
  NAND2_X1 U73 ( .A1(n113), .A2(n112), .ZN(C[23]) );
  INV_X1 U74 ( .A(B[24]), .ZN(n114) );
  NAND2_X1 U75 ( .A1(n114), .A2(n86), .ZN(C[24]) );
  INV_X1 U76 ( .A(B[25]), .ZN(n115) );
  NAND2_X1 U77 ( .A1(n115), .A2(n87), .ZN(C[25]) );
  INV_X1 U78 ( .A(B[26]), .ZN(n116) );
  NAND2_X1 U79 ( .A1(n116), .A2(n88), .ZN(C[26]) );
  INV_X1 U80 ( .A(B[27]), .ZN(n118) );
  INV_X1 U81 ( .A(A[27]), .ZN(n117) );
  NAND2_X1 U82 ( .A1(n118), .A2(n117), .ZN(C[27]) );
  INV_X1 U83 ( .A(B[28]), .ZN(n120) );
  INV_X1 U84 ( .A(A[28]), .ZN(n119) );
  NAND2_X1 U85 ( .A1(n120), .A2(n119), .ZN(C[28]) );
  INV_X1 U86 ( .A(B[29]), .ZN(n122) );
  INV_X1 U87 ( .A(A[29]), .ZN(n121) );
  NAND2_X1 U88 ( .A1(n122), .A2(n121), .ZN(C[29]) );
  INV_X1 U89 ( .A(B[30]), .ZN(n124) );
  INV_X1 U90 ( .A(A[30]), .ZN(n123) );
  NAND2_X1 U91 ( .A1(n124), .A2(n123), .ZN(C[30]) );
  INV_X1 U92 ( .A(B[31]), .ZN(n126) );
  INV_X1 U93 ( .A(A[31]), .ZN(n125) );
  NAND2_X1 U94 ( .A1(n126), .A2(n125), .ZN(C[31]) );
endmodule


module and_gen_N32 ( A, B, C );
  input [31:0] A;
  input [31:0] B;
  output [31:0] C;


  AND2_X1 U1 ( .A1(A[15]), .A2(B[15]), .ZN(C[15]) );
  AND2_X1 U2 ( .A1(A[1]), .A2(B[1]), .ZN(C[1]) );
  AND2_X1 U3 ( .A1(A[23]), .A2(B[23]), .ZN(C[23]) );
  AND2_X1 U4 ( .A1(A[21]), .A2(B[21]), .ZN(C[21]) );
  AND2_X1 U5 ( .A1(A[17]), .A2(B[17]), .ZN(C[17]) );
  AND2_X1 U6 ( .A1(A[28]), .A2(B[28]), .ZN(C[28]) );
  AND2_X1 U7 ( .A1(A[16]), .A2(B[16]), .ZN(C[16]) );
  AND2_X1 U8 ( .A1(A[19]), .A2(B[19]), .ZN(C[19]) );
  AND2_X1 U9 ( .A1(A[27]), .A2(B[27]), .ZN(C[27]) );
  AND2_X1 U10 ( .A1(A[29]), .A2(B[29]), .ZN(C[29]) );
  AND2_X1 U11 ( .A1(A[18]), .A2(B[18]), .ZN(C[18]) );
  AND2_X1 U12 ( .A1(A[30]), .A2(B[30]), .ZN(C[30]) );
  AND2_X1 U13 ( .A1(A[2]), .A2(B[2]), .ZN(C[2]) );
  AND2_X1 U14 ( .A1(A[31]), .A2(B[31]), .ZN(C[31]) );
  AND2_X1 U15 ( .A1(A[22]), .A2(B[22]), .ZN(C[22]) );
  AND2_X1 U16 ( .A1(A[14]), .A2(B[14]), .ZN(C[14]) );
  AND2_X1 U17 ( .A1(A[13]), .A2(B[13]), .ZN(C[13]) );
  AND2_X1 U18 ( .A1(A[24]), .A2(B[24]), .ZN(C[24]) );
  AND2_X1 U19 ( .A1(A[25]), .A2(B[25]), .ZN(C[25]) );
  AND2_X1 U20 ( .A1(A[26]), .A2(B[26]), .ZN(C[26]) );
  AND2_X1 U21 ( .A1(A[3]), .A2(B[3]), .ZN(C[3]) );
  AND2_X1 U22 ( .A1(A[20]), .A2(B[20]), .ZN(C[20]) );
  AND2_X1 U23 ( .A1(A[11]), .A2(B[11]), .ZN(C[11]) );
  AND2_X1 U24 ( .A1(A[12]), .A2(B[12]), .ZN(C[12]) );
  AND2_X1 U25 ( .A1(A[10]), .A2(B[10]), .ZN(C[10]) );
  AND2_X1 U26 ( .A1(A[5]), .A2(B[5]), .ZN(C[5]) );
  AND2_X1 U27 ( .A1(A[7]), .A2(B[7]), .ZN(C[7]) );
  AND2_X1 U28 ( .A1(A[4]), .A2(B[4]), .ZN(C[4]) );
  AND2_X1 U29 ( .A1(A[8]), .A2(B[8]), .ZN(C[8]) );
  AND2_X1 U30 ( .A1(A[0]), .A2(B[0]), .ZN(C[0]) );
  AND2_X1 U31 ( .A1(A[6]), .A2(B[6]), .ZN(C[6]) );
  AND2_X1 U32 ( .A1(A[9]), .A2(B[9]), .ZN(C[9]) );
endmodule


module MUX21_GENERIC_N32_12 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_647 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n6), .Y(Y[0]) );
  MUX21_646 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n5), .Y(Y[1]) );
  MUX21_645 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_644 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n6), .Y(Y[3]) );
  MUX21_643 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n6), .Y(Y[4]) );
  MUX21_642 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n6), .Y(Y[5]) );
  MUX21_641 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_640 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n6), .Y(Y[7]) );
  MUX21_639 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_638 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n6), .Y(Y[9]) );
  MUX21_637 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_636 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n6), .Y(Y[11]) );
  MUX21_635 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n4), .Y(Y[12]) );
  MUX21_634 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n6), .Y(Y[13]) );
  MUX21_633 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n4), .Y(Y[14]) );
  MUX21_632 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n4), .Y(Y[15]) );
  MUX21_631 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n4), .Y(Y[16]) );
  MUX21_630 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n4), .Y(Y[17]) );
  MUX21_629 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n4), .Y(Y[18]) );
  MUX21_628 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n4), .Y(Y[19]) );
  MUX21_627 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n4), .Y(Y[20]) );
  MUX21_626 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_625 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_624 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_623 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n5), .Y(Y[24]) );
  MUX21_622 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n5), .Y(Y[25]) );
  MUX21_621 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n5), .Y(Y[26]) );
  MUX21_620 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n5), .Y(Y[27]) );
  MUX21_619 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n5), .Y(Y[28]) );
  MUX21_618 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n5), .Y(Y[29]) );
  MUX21_617 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n5), .Y(Y[30]) );
  MUX21_616 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n5), .Y(Y[31]) );
  BUF_X2 U1 ( .A(n3), .Z(n6) );
  BUF_X4 U2 ( .A(n3), .Z(n4) );
  BUF_X4 U3 ( .A(n3), .Z(n5) );
endmodule


module MUX21_GENERIC_N32_13 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n2, n3, n4, n5, n6;
  assign n2 = S;

  MUX21_679 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_678 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_677 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_676 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_675 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n5), .Y(Y[4]) );
  MUX21_674 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n6), .Y(Y[5]) );
  MUX21_673 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n5), .Y(Y[6]) );
  MUX21_672 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n3), .Y(Y[7]) );
  MUX21_671 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n5), .Y(Y[8]) );
  MUX21_670 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n6), .Y(Y[9]) );
  MUX21_669 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n5), .Y(Y[10]) );
  MUX21_668 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n3), .Y(Y[11]) );
  MUX21_667 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_666 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n6), .Y(Y[13]) );
  MUX21_665 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_664 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n3), .Y(Y[15]) );
  MUX21_663 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_662 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n6), .Y(Y[17]) );
  MUX21_661 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n3), .Y(Y[18]) );
  MUX21_660 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_659 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_658 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n6), .Y(Y[21]) );
  MUX21_657 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_656 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_655 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_654 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_653 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n5), .Y(Y[26]) );
  MUX21_652 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_651 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_650 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_649 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_648 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(n5), .Z(n6) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n3) );
  BUF_X2 U3 ( .A(n2), .Z(n4) );
  BUF_X4 U4 ( .A(n2), .Z(n5) );
endmodule


module MUX21_GENERIC_N32_14 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5;
  assign n3 = S;

  MUX21_711 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_710 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_709 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_708 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_707 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n5), .Y(Y[4]) );
  MUX21_706 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n5), .Y(Y[5]) );
  MUX21_705 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n5), .Y(Y[6]) );
  MUX21_704 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n5), .Y(Y[7]) );
  MUX21_703 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n5), .Y(Y[8]) );
  MUX21_702 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n5), .Y(Y[9]) );
  MUX21_701 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n5), .Y(Y[10]) );
  MUX21_700 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n5), .Y(Y[11]) );
  MUX21_699 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_698 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_697 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_696 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_695 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_694 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_693 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_692 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_691 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_690 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_689 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_688 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_687 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n5), .Y(Y[24]) );
  MUX21_686 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n5), .Y(Y[25]) );
  MUX21_685 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n5), .Y(Y[26]) );
  MUX21_684 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n5), .Y(Y[27]) );
  MUX21_683 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n5), .Y(Y[28]) );
  MUX21_682 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n5), .Y(Y[29]) );
  MUX21_681 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n5), .Y(Y[30]) );
  MUX21_680 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n5), .Y(Y[31]) );
  BUF_X2 U1 ( .A(n3), .Z(n4) );
  BUF_X8 U2 ( .A(n3), .Z(n5) );
endmodule


module MUX21_GENERIC_N32_15 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_743 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n6), .Y(Y[0]) );
  MUX21_742 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n6), .Y(Y[1]) );
  MUX21_741 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n5), .Y(Y[2]) );
  MUX21_740 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n5), .Y(Y[3]) );
  MUX21_739 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n5), .Y(Y[4]) );
  MUX21_738 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_737 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_736 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_735 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n5), .Y(Y[8]) );
  MUX21_734 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_733 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_732 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n5), .Y(Y[11]) );
  MUX21_731 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n4), .Y(Y[12]) );
  MUX21_730 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n4), .Y(Y[13]) );
  MUX21_729 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n6), .Y(Y[14]) );
  MUX21_728 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n4), .Y(Y[15]) );
  MUX21_727 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n4), .Y(Y[16]) );
  MUX21_726 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n4), .Y(Y[17]) );
  MUX21_725 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n6), .Y(Y[18]) );
  MUX21_724 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n6), .Y(Y[19]) );
  MUX21_723 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n4), .Y(Y[20]) );
  MUX21_722 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n4), .Y(Y[21]) );
  MUX21_721 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_720 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_719 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n5), .Y(Y[24]) );
  MUX21_718 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n5), .Y(Y[25]) );
  MUX21_717 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n5), .Y(Y[26]) );
  MUX21_716 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n5), .Y(Y[27]) );
  MUX21_715 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_714 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_713 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_712 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n5), .Y(Y[31]) );
  BUF_X2 U1 ( .A(n3), .Z(n6) );
  BUF_X4 U2 ( .A(n3), .Z(n4) );
  BUF_X4 U3 ( .A(n3), .Z(n5) );
endmodule


module MUX21_GENERIC_N32_16 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n7, n8, n9, n10, n11, n12;
  assign n7 = S;

  MUX21_775 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n8), .Y(Y[0]) );
  MUX21_774 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n12), .Y(Y[1]) );
  MUX21_773 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n12), .Y(Y[2]) );
  MUX21_772 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n12), .Y(Y[3]) );
  MUX21_771 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n10), .Y(Y[4]) );
  MUX21_770 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n12), .Y(Y[5]) );
  MUX21_769 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n8), .Y(Y[6]) );
  MUX21_768 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n10), .Y(Y[7]) );
  MUX21_767 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n8), .Y(Y[8]) );
  MUX21_766 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n10), .Y(Y[9]) );
  MUX21_765 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n8), .Y(Y[10]) );
  MUX21_764 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n10), .Y(Y[11]) );
  MUX21_763 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n10), .Y(Y[12]) );
  MUX21_762 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n9), .Y(Y[13]) );
  MUX21_761 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n11), .Y(Y[14]) );
  MUX21_760 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n11), .Y(Y[15]) );
  MUX21_759 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n11), .Y(Y[16]) );
  MUX21_758 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n11), .Y(Y[17]) );
  MUX21_757 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n11), .Y(Y[18]) );
  MUX21_756 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n11), .Y(Y[19]) );
  MUX21_755 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n11), .Y(Y[20]) );
  MUX21_754 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n11), .Y(Y[21]) );
  MUX21_753 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n11), .Y(Y[22]) );
  MUX21_752 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n11), .Y(Y[23]) );
  MUX21_751 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n11), .Y(Y[24]) );
  MUX21_750 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n11), .Y(Y[25]) );
  MUX21_749 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n12), .Y(Y[26]) );
  MUX21_748 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n10), .Y(Y[27]) );
  MUX21_747 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n11), .Y(Y[28]) );
  MUX21_746 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n8), .Y(Y[29]) );
  MUX21_745 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n11), .Y(Y[30]) );
  MUX21_744 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n11), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(n7), .Z(n12) );
  CLKBUF_X3 U2 ( .A(n7), .Z(n10) );
  CLKBUF_X3 U3 ( .A(n7), .Z(n8) );
  BUF_X4 U4 ( .A(n8), .Z(n11) );
  BUF_X1 U5 ( .A(n12), .Z(n9) );
endmodule


module MUX21_GENERIC_N32_17 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n5, n6, n7, n8;
  assign n5 = S;

  MUX21_807 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n7), .Y(Y[0]) );
  MUX21_806 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n7), .Y(Y[1]) );
  MUX21_805 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n8), .Y(Y[2]) );
  MUX21_804 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n7), .Y(Y[3]) );
  MUX21_803 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n6), .Y(Y[4]) );
  MUX21_802 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n8), .Y(Y[5]) );
  MUX21_801 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n7), .Y(Y[6]) );
  MUX21_800 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n7), .Y(Y[7]) );
  MUX21_799 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n8), .Y(Y[8]) );
  MUX21_798 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n7), .Y(Y[9]) );
  MUX21_797 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n8), .Y(Y[10]) );
  MUX21_796 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n6), .Y(Y[11]) );
  MUX21_795 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n6), .Y(Y[12]) );
  MUX21_794 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n6), .Y(Y[13]) );
  MUX21_793 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n8), .Y(Y[14]) );
  MUX21_792 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n6), .Y(Y[15]) );
  MUX21_791 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n6), .Y(Y[16]) );
  MUX21_790 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n8), .Y(Y[17]) );
  MUX21_789 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n8), .Y(Y[18]) );
  MUX21_788 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n8), .Y(Y[19]) );
  MUX21_787 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n8), .Y(Y[20]) );
  MUX21_786 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n6), .Y(Y[21]) );
  MUX21_785 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n6), .Y(Y[22]) );
  MUX21_784 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n6), .Y(Y[23]) );
  MUX21_783 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n8), .Y(Y[24]) );
  MUX21_782 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n8), .Y(Y[25]) );
  MUX21_781 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_780 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_779 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_778 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n8), .Y(Y[29]) );
  MUX21_777 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_776 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n8), .Y(Y[31]) );
  CLKBUF_X3 U1 ( .A(n5), .Z(n7) );
  BUF_X4 U2 ( .A(n5), .Z(n6) );
  BUF_X4 U3 ( .A(n5), .Z(n8) );
endmodule


module MUX21_GENERIC_N32_18 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_839 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_838 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_837 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_836 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_835 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_834 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_833 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_832 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_831 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_830 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_829 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_828 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_827 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_826 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_825 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_824 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_823 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n5), .Y(Y[16]) );
  MUX21_822 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_821 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_820 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_819 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_818 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_817 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_816 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_815 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n6), .Y(Y[24]) );
  MUX21_814 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_813 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_812 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_811 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_810 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_809 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_808 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n5) );
  BUF_X1 U2 ( .A(n3), .Z(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_19 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_871 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n5), .Y(Y[0]) );
  MUX21_870 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n5), .Y(Y[1]) );
  MUX21_869 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n5), .Y(Y[2]) );
  MUX21_868 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n5), .Y(Y[3]) );
  MUX21_867 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n5), .Y(Y[4]) );
  MUX21_866 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n5), .Y(Y[5]) );
  MUX21_865 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n5), .Y(Y[6]) );
  MUX21_864 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n5), .Y(Y[7]) );
  MUX21_863 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n6), .Y(Y[8]) );
  MUX21_862 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n6), .Y(Y[9]) );
  MUX21_861 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n6), .Y(Y[10]) );
  MUX21_860 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n6), .Y(Y[11]) );
  MUX21_859 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n6), .Y(Y[12]) );
  MUX21_858 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n6), .Y(Y[13]) );
  MUX21_857 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n6), .Y(Y[14]) );
  MUX21_856 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n6), .Y(Y[15]) );
  MUX21_855 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n4), .Y(Y[16]) );
  MUX21_854 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n4), .Y(Y[17]) );
  MUX21_853 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n4), .Y(Y[18]) );
  MUX21_852 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n4), .Y(Y[19]) );
  MUX21_851 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n4), .Y(Y[20]) );
  MUX21_850 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n4), .Y(Y[21]) );
  MUX21_849 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n4), .Y(Y[22]) );
  MUX21_848 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n4), .Y(Y[23]) );
  MUX21_847 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n4), .Y(Y[24]) );
  MUX21_846 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n4), .Y(Y[25]) );
  MUX21_845 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n4), .Y(Y[26]) );
  MUX21_844 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n4), .Y(Y[27]) );
  MUX21_843 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n5), .Y(Y[28]) );
  MUX21_842 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n5), .Y(Y[29]) );
  MUX21_841 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n5), .Y(Y[30]) );
  MUX21_840 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n5), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n5) );
  BUF_X1 U2 ( .A(n3), .Z(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module MUX21_GENERIC_N32_0 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   n3, n4, n5, n6;
  assign n3 = S;

  MUX21_903 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n4), .Y(Y[0]) );
  MUX21_902 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n4), .Y(Y[1]) );
  MUX21_901 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n4), .Y(Y[2]) );
  MUX21_900 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n4), .Y(Y[3]) );
  MUX21_899 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n4), .Y(Y[4]) );
  MUX21_898 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n4), .Y(Y[5]) );
  MUX21_897 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n4), .Y(Y[6]) );
  MUX21_896 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n4), .Y(Y[7]) );
  MUX21_895 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n4), .Y(Y[8]) );
  MUX21_894 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n4), .Y(Y[9]) );
  MUX21_893 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n4), .Y(Y[10]) );
  MUX21_892 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n4), .Y(Y[11]) );
  MUX21_891 MUXes_12 ( .A(A[12]), .B(B[12]), .S(n5), .Y(Y[12]) );
  MUX21_890 MUXes_13 ( .A(A[13]), .B(B[13]), .S(n5), .Y(Y[13]) );
  MUX21_889 MUXes_14 ( .A(A[14]), .B(B[14]), .S(n5), .Y(Y[14]) );
  MUX21_888 MUXes_15 ( .A(A[15]), .B(B[15]), .S(n5), .Y(Y[15]) );
  MUX21_887 MUXes_16 ( .A(A[16]), .B(B[16]), .S(n6), .Y(Y[16]) );
  MUX21_886 MUXes_17 ( .A(A[17]), .B(B[17]), .S(n5), .Y(Y[17]) );
  MUX21_885 MUXes_18 ( .A(A[18]), .B(B[18]), .S(n5), .Y(Y[18]) );
  MUX21_884 MUXes_19 ( .A(A[19]), .B(B[19]), .S(n5), .Y(Y[19]) );
  MUX21_883 MUXes_20 ( .A(A[20]), .B(B[20]), .S(n5), .Y(Y[20]) );
  MUX21_882 MUXes_21 ( .A(A[21]), .B(B[21]), .S(n5), .Y(Y[21]) );
  MUX21_881 MUXes_22 ( .A(A[22]), .B(B[22]), .S(n5), .Y(Y[22]) );
  MUX21_880 MUXes_23 ( .A(A[23]), .B(B[23]), .S(n5), .Y(Y[23]) );
  MUX21_879 MUXes_24 ( .A(A[24]), .B(B[24]), .S(n5), .Y(Y[24]) );
  MUX21_878 MUXes_25 ( .A(A[25]), .B(B[25]), .S(n6), .Y(Y[25]) );
  MUX21_877 MUXes_26 ( .A(A[26]), .B(B[26]), .S(n6), .Y(Y[26]) );
  MUX21_876 MUXes_27 ( .A(A[27]), .B(B[27]), .S(n6), .Y(Y[27]) );
  MUX21_875 MUXes_28 ( .A(A[28]), .B(B[28]), .S(n6), .Y(Y[28]) );
  MUX21_874 MUXes_29 ( .A(A[29]), .B(B[29]), .S(n6), .Y(Y[29]) );
  MUX21_873 MUXes_30 ( .A(A[30]), .B(B[30]), .S(n6), .Y(Y[30]) );
  MUX21_872 MUXes_31 ( .A(A[31]), .B(B[31]), .S(n6), .Y(Y[31]) );
  BUF_X1 U1 ( .A(n3), .Z(n5) );
  BUF_X1 U2 ( .A(n3), .Z(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n6) );
endmodule


module MUX21_GENERIC_N5_1 ( A, B, S, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input S;


  MUX21_908 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_907 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_906 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_905 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
  MUX21_904 MUXes_4 ( .A(A[4]), .B(B[4]), .S(S), .Y(Y[4]) );
endmodule


module MUX21_GENERIC_N5_2 ( A, B, S, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input S;


  MUX21_913 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_912 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_911 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_910 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
  MUX21_909 MUXes_4 ( .A(A[4]), .B(B[4]), .S(S), .Y(Y[4]) );
endmodule


module MUX21_GENERIC_N5_0 ( A, B, S, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input S;


  MUX21_918 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_917 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_916 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_915 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
  MUX21_914 MUXes_4 ( .A(A[4]), .B(B[4]), .S(S), .Y(Y[4]) );
endmodule


module FA_523 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n8, n9, n10, n11;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n11) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n10) );
  INV_X1 U3 ( .A(n11), .ZN(n8) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n10), .A2(n9), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n11), .ZN(S) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n7, n8, n9;

  XOR2_X1 U1 ( .A(n8), .B(n9), .Z(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n8) );
  OAI21_X1 U3 ( .B1(n8), .B2(n9), .A(n7), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n9) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
endmodule


module MUX21_921 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_921 UIV ( .A(S), .Y(SB) );
  ND2_2763 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2762 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2761 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_931 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_931 UIV ( .A(S), .Y(SB) );
  ND2_2793 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2792 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2791 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_942 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_942 UIV ( .A(S), .Y(SB) );
  ND2_2826 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2825 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2824 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   SB, Y1, Y2;

  IV_0 UIV ( .A(S), .Y(SB) );
  ND2_0 UND1 ( .A(A), .B(SB), .Y(Y1) );
  ND2_2828 UND2 ( .A(B), .B(S), .Y(Y2) );
  ND2_2827 UND3 ( .A(Y1), .B(Y2), .Y(Y) );
endmodule


module mux41_generic_N32_1 ( A, B, C, D, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Y;

  wire   [31:0] ABto2;
  wire   [31:0] CDto2;

  MUX21_GENERIC_N32_10 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_GENERIC_N32_9 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_GENERIC_N32_8 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(Y) );
endmodule


module D_Reg_generic_N5_1 ( D, CLK, RESET, ENABLE, Q );
  input [4:0] D;
  output [4:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, net56157, net56158, net56159, net56160, net56161,
         n6, n7, n8, n9, n10, n17;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(CLK), .RN(RESET), .Q(Q[4]), .QN(net56161)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(CLK), .RN(RESET), .Q(Q[3]), .QN(net56160)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(CLK), .RN(RESET), .Q(Q[2]), .QN(net56159)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(CLK), .RN(RESET), .Q(Q[1]), .QN(net56158)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(CLK), .RN(RESET), .Q(Q[0]), .QN(net56157)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n17) );
  OAI21_X1 U3 ( .B1(net56157), .B2(n17), .A(n6), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n17), .A2(D[0]), .ZN(n6) );
  OAI21_X1 U5 ( .B1(net56158), .B2(n17), .A(n7), .ZN(n4) );
  NAND2_X1 U6 ( .A1(D[1]), .A2(n17), .ZN(n7) );
  OAI21_X1 U7 ( .B1(net56159), .B2(n17), .A(n8), .ZN(n3) );
  NAND2_X1 U8 ( .A1(D[2]), .A2(n17), .ZN(n8) );
  OAI21_X1 U9 ( .B1(net56160), .B2(n17), .A(n9), .ZN(n2) );
  NAND2_X1 U10 ( .A1(D[3]), .A2(n17), .ZN(n9) );
  OAI21_X1 U11 ( .B1(net56161), .B2(n17), .A(n10), .ZN(n1) );
  NAND2_X1 U12 ( .A1(D[4]), .A2(n17), .ZN(n10) );
endmodule


module D_Reg_generic_N32_1 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55837, net55838, net55839, net55840, net55841, net55842,
         net55843, net55844, net55845, net55846, net55847, net55848, net55849,
         net55850, net55851, net55852, net55853, net55854, net55855, net55856,
         net55857, net55858, net55859, net55860, net55861, net55862, net55863,
         net55864, net55865, net55866, net55867, net55868, n73, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n106, n107, n108, n109, n110, n111, n112, n113, n114;
  assign n73 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n114), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n112), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n114), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n112), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n114), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n112), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n112), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n112), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n114), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n112), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n112), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n112), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n114), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n113), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n113), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n113), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n112), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n113), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n113), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n113), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n113), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n113), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n114), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n112), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n114), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n112), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n113), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n112), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n113), .Q(Q[3]), .QN(net55840)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n113), .Q(Q[2]), .QN(net55839)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n113), .Q(Q[1]), .QN(net55838)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n114), .Q(Q[0]), .QN(net55837)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n106) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n107) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n108) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n110) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n109) );
  OAI21_X1 U7 ( .B1(net55860), .B2(n109), .A(n33), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n111), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U9 ( .B1(net55845), .B2(n109), .A(n48), .ZN(n24) );
  NAND2_X1 U10 ( .A1(D[8]), .A2(n108), .ZN(n48) );
  OAI21_X1 U11 ( .B1(net55846), .B2(n110), .A(n49), .ZN(n23) );
  NAND2_X1 U12 ( .A1(D[9]), .A2(n108), .ZN(n49) );
  OAI21_X1 U13 ( .B1(net55868), .B2(n109), .A(n64), .ZN(n1) );
  NAND2_X1 U14 ( .A1(D[31]), .A2(n106), .ZN(n64) );
  OAI21_X1 U15 ( .B1(net55837), .B2(n109), .A(n39), .ZN(n32) );
  NAND2_X1 U16 ( .A1(D[0]), .A2(n107), .ZN(n39) );
  OAI21_X1 U17 ( .B1(net55838), .B2(n108), .A(n40), .ZN(n31) );
  NAND2_X1 U18 ( .A1(D[1]), .A2(n107), .ZN(n40) );
  OAI21_X1 U19 ( .B1(net55839), .B2(n109), .A(n41), .ZN(n30) );
  NAND2_X1 U20 ( .A1(D[2]), .A2(n107), .ZN(n41) );
  OAI21_X1 U21 ( .B1(net55840), .B2(n109), .A(n43), .ZN(n29) );
  NAND2_X1 U22 ( .A1(D[3]), .A2(n107), .ZN(n43) );
  OAI21_X1 U23 ( .B1(net55857), .B2(n111), .A(n61), .ZN(n12) );
  NAND2_X1 U24 ( .A1(D[20]), .A2(n106), .ZN(n61) );
  OAI21_X1 U25 ( .B1(net55858), .B2(n111), .A(n62), .ZN(n11) );
  NAND2_X1 U26 ( .A1(D[21]), .A2(n106), .ZN(n62) );
  OAI21_X1 U27 ( .B1(net55859), .B2(n111), .A(n63), .ZN(n10) );
  NAND2_X1 U28 ( .A1(D[22]), .A2(n106), .ZN(n63) );
  OAI21_X1 U29 ( .B1(net55847), .B2(n110), .A(n50), .ZN(n22) );
  NAND2_X1 U30 ( .A1(D[10]), .A2(n107), .ZN(n50) );
  OAI21_X1 U31 ( .B1(net55848), .B2(n110), .A(n51), .ZN(n21) );
  NAND2_X1 U32 ( .A1(D[11]), .A2(n107), .ZN(n51) );
  OAI21_X1 U33 ( .B1(net55849), .B2(n110), .A(n52), .ZN(n20) );
  NAND2_X1 U34 ( .A1(D[12]), .A2(n107), .ZN(n52) );
  OAI21_X1 U35 ( .B1(net55850), .B2(n110), .A(n54), .ZN(n19) );
  NAND2_X1 U36 ( .A1(D[13]), .A2(n107), .ZN(n54) );
  OAI21_X1 U37 ( .B1(net55851), .B2(n110), .A(n55), .ZN(n18) );
  NAND2_X1 U38 ( .A1(D[14]), .A2(n107), .ZN(n55) );
  OAI21_X1 U39 ( .B1(net55852), .B2(n110), .A(n56), .ZN(n17) );
  NAND2_X1 U40 ( .A1(D[15]), .A2(n107), .ZN(n56) );
  OAI21_X1 U41 ( .B1(net55853), .B2(n110), .A(n57), .ZN(n16) );
  NAND2_X1 U42 ( .A1(D[16]), .A2(n106), .ZN(n57) );
  OAI21_X1 U43 ( .B1(net55854), .B2(n110), .A(n58), .ZN(n15) );
  NAND2_X1 U44 ( .A1(D[17]), .A2(n106), .ZN(n58) );
  OAI21_X1 U45 ( .B1(net55855), .B2(n110), .A(n59), .ZN(n14) );
  NAND2_X1 U46 ( .A1(D[18]), .A2(n106), .ZN(n59) );
  OAI21_X1 U47 ( .B1(net55856), .B2(n110), .A(n60), .ZN(n13) );
  NAND2_X1 U48 ( .A1(D[19]), .A2(n106), .ZN(n60) );
  OAI21_X1 U49 ( .B1(net55861), .B2(n108), .A(n34), .ZN(n8) );
  NAND2_X1 U50 ( .A1(D[24]), .A2(n106), .ZN(n34) );
  OAI21_X1 U51 ( .B1(net55862), .B2(n108), .A(n35), .ZN(n7) );
  NAND2_X1 U52 ( .A1(D[25]), .A2(n106), .ZN(n35) );
  OAI21_X1 U53 ( .B1(net55863), .B2(n109), .A(n36), .ZN(n6) );
  NAND2_X1 U54 ( .A1(D[26]), .A2(n106), .ZN(n36) );
  OAI21_X1 U55 ( .B1(net55864), .B2(n108), .A(n37), .ZN(n5) );
  NAND2_X1 U56 ( .A1(D[27]), .A2(n106), .ZN(n37) );
  OAI21_X1 U57 ( .B1(net55865), .B2(n108), .A(n38), .ZN(n4) );
  NAND2_X1 U58 ( .A1(D[28]), .A2(n107), .ZN(n38) );
  OAI21_X1 U59 ( .B1(net55867), .B2(n110), .A(n53), .ZN(n2) );
  NAND2_X1 U60 ( .A1(D[30]), .A2(n107), .ZN(n53) );
  OAI21_X1 U61 ( .B1(net55841), .B2(n109), .A(n44), .ZN(n28) );
  NAND2_X1 U62 ( .A1(D[4]), .A2(n108), .ZN(n44) );
  OAI21_X1 U63 ( .B1(net55842), .B2(n109), .A(n45), .ZN(n27) );
  NAND2_X1 U64 ( .A1(D[5]), .A2(n108), .ZN(n45) );
  OAI21_X1 U65 ( .B1(net55843), .B2(n109), .A(n46), .ZN(n26) );
  NAND2_X1 U66 ( .A1(D[6]), .A2(n108), .ZN(n46) );
  OAI21_X1 U67 ( .B1(net55844), .B2(n109), .A(n47), .ZN(n25) );
  NAND2_X1 U68 ( .A1(D[7]), .A2(n108), .ZN(n47) );
  OAI21_X1 U69 ( .B1(net55866), .B2(n109), .A(n42), .ZN(n3) );
  NAND2_X1 U70 ( .A1(D[29]), .A2(n108), .ZN(n42) );
  BUF_X1 U71 ( .A(n73), .Z(n113) );
  BUF_X1 U72 ( .A(n73), .Z(n112) );
  BUF_X1 U73 ( .A(n73), .Z(n114) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n111) );
endmodule


module D_Reg_generic_N32_2 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55837, net55838, net55839, net55840, net55841, net55842,
         net55843, net55844, net55845, net55846, net55847, net55848, net55849,
         net55850, net55851, net55852, net55853, net55854, net55855, net55856,
         net55857, net55858, net55859, net55860, net55861, net55862, net55863,
         net55864, net55865, net55866, net55867, net55868, n73, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n106, n107, n108, n109, n110, n111, n112, n113, n114;
  assign n73 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n114), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n112), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n114), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n112), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n114), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n112), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n112), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n112), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n114), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n112), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n112), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n112), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n114), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n113), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n113), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n113), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n112), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n113), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n113), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n113), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n113), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n113), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n114), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n112), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n114), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n112), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n113), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n112), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n113), .Q(Q[3]), .QN(net55840)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n113), .Q(Q[2]), .QN(net55839)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n113), .Q(Q[1]), .QN(net55838)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n114), .Q(Q[0]), .QN(net55837)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n106) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n107) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n108) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n110) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n109) );
  OAI21_X1 U7 ( .B1(net55860), .B2(n109), .A(n33), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n111), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U9 ( .B1(net55841), .B2(n109), .A(n44), .ZN(n28) );
  NAND2_X1 U10 ( .A1(D[4]), .A2(n108), .ZN(n44) );
  OAI21_X1 U11 ( .B1(net55842), .B2(n109), .A(n45), .ZN(n27) );
  NAND2_X1 U12 ( .A1(D[5]), .A2(n108), .ZN(n45) );
  OAI21_X1 U13 ( .B1(net55843), .B2(n109), .A(n46), .ZN(n26) );
  NAND2_X1 U14 ( .A1(D[6]), .A2(n108), .ZN(n46) );
  OAI21_X1 U15 ( .B1(net55844), .B2(n109), .A(n47), .ZN(n25) );
  NAND2_X1 U16 ( .A1(D[7]), .A2(n108), .ZN(n47) );
  OAI21_X1 U17 ( .B1(net55845), .B2(n109), .A(n48), .ZN(n24) );
  NAND2_X1 U18 ( .A1(D[8]), .A2(n108), .ZN(n48) );
  OAI21_X1 U19 ( .B1(net55846), .B2(n110), .A(n49), .ZN(n23) );
  NAND2_X1 U20 ( .A1(D[9]), .A2(n108), .ZN(n49) );
  OAI21_X1 U21 ( .B1(net55866), .B2(n109), .A(n42), .ZN(n3) );
  NAND2_X1 U22 ( .A1(D[29]), .A2(n108), .ZN(n42) );
  OAI21_X1 U23 ( .B1(net55857), .B2(n111), .A(n61), .ZN(n12) );
  NAND2_X1 U24 ( .A1(D[20]), .A2(n106), .ZN(n61) );
  OAI21_X1 U25 ( .B1(net55858), .B2(n111), .A(n62), .ZN(n11) );
  NAND2_X1 U26 ( .A1(D[21]), .A2(n106), .ZN(n62) );
  OAI21_X1 U27 ( .B1(net55859), .B2(n111), .A(n63), .ZN(n10) );
  NAND2_X1 U28 ( .A1(D[22]), .A2(n106), .ZN(n63) );
  OAI21_X1 U29 ( .B1(net55838), .B2(n108), .A(n40), .ZN(n31) );
  NAND2_X1 U30 ( .A1(D[1]), .A2(n107), .ZN(n40) );
  OAI21_X1 U31 ( .B1(net55861), .B2(n108), .A(n34), .ZN(n8) );
  NAND2_X1 U32 ( .A1(D[24]), .A2(n106), .ZN(n34) );
  OAI21_X1 U33 ( .B1(net55862), .B2(n108), .A(n35), .ZN(n7) );
  NAND2_X1 U34 ( .A1(D[25]), .A2(n106), .ZN(n35) );
  OAI21_X1 U35 ( .B1(net55864), .B2(n108), .A(n37), .ZN(n5) );
  NAND2_X1 U36 ( .A1(D[27]), .A2(n106), .ZN(n37) );
  OAI21_X1 U37 ( .B1(net55865), .B2(n108), .A(n38), .ZN(n4) );
  NAND2_X1 U38 ( .A1(D[28]), .A2(n107), .ZN(n38) );
  OAI21_X1 U39 ( .B1(net55837), .B2(n109), .A(n39), .ZN(n32) );
  NAND2_X1 U40 ( .A1(D[0]), .A2(n107), .ZN(n39) );
  OAI21_X1 U41 ( .B1(net55839), .B2(n109), .A(n41), .ZN(n30) );
  NAND2_X1 U42 ( .A1(D[2]), .A2(n107), .ZN(n41) );
  OAI21_X1 U43 ( .B1(net55840), .B2(n109), .A(n43), .ZN(n29) );
  NAND2_X1 U44 ( .A1(D[3]), .A2(n107), .ZN(n43) );
  OAI21_X1 U45 ( .B1(net55847), .B2(n110), .A(n50), .ZN(n22) );
  NAND2_X1 U46 ( .A1(D[10]), .A2(n107), .ZN(n50) );
  OAI21_X1 U47 ( .B1(net55848), .B2(n110), .A(n51), .ZN(n21) );
  NAND2_X1 U48 ( .A1(D[11]), .A2(n107), .ZN(n51) );
  OAI21_X1 U49 ( .B1(net55849), .B2(n110), .A(n52), .ZN(n20) );
  NAND2_X1 U50 ( .A1(D[12]), .A2(n107), .ZN(n52) );
  OAI21_X1 U51 ( .B1(net55850), .B2(n110), .A(n54), .ZN(n19) );
  NAND2_X1 U52 ( .A1(D[13]), .A2(n107), .ZN(n54) );
  OAI21_X1 U53 ( .B1(net55851), .B2(n110), .A(n55), .ZN(n18) );
  NAND2_X1 U54 ( .A1(D[14]), .A2(n107), .ZN(n55) );
  OAI21_X1 U55 ( .B1(net55852), .B2(n110), .A(n56), .ZN(n17) );
  NAND2_X1 U56 ( .A1(D[15]), .A2(n107), .ZN(n56) );
  OAI21_X1 U57 ( .B1(net55853), .B2(n110), .A(n57), .ZN(n16) );
  NAND2_X1 U58 ( .A1(D[16]), .A2(n106), .ZN(n57) );
  OAI21_X1 U59 ( .B1(net55854), .B2(n110), .A(n58), .ZN(n15) );
  NAND2_X1 U60 ( .A1(D[17]), .A2(n106), .ZN(n58) );
  OAI21_X1 U61 ( .B1(net55855), .B2(n110), .A(n59), .ZN(n14) );
  NAND2_X1 U62 ( .A1(D[18]), .A2(n106), .ZN(n59) );
  OAI21_X1 U63 ( .B1(net55856), .B2(n110), .A(n60), .ZN(n13) );
  NAND2_X1 U64 ( .A1(D[19]), .A2(n106), .ZN(n60) );
  OAI21_X1 U65 ( .B1(net55863), .B2(n109), .A(n36), .ZN(n6) );
  NAND2_X1 U66 ( .A1(D[26]), .A2(n106), .ZN(n36) );
  OAI21_X1 U67 ( .B1(net55867), .B2(n110), .A(n53), .ZN(n2) );
  NAND2_X1 U68 ( .A1(D[30]), .A2(n107), .ZN(n53) );
  OAI21_X1 U69 ( .B1(net55868), .B2(n109), .A(n64), .ZN(n1) );
  NAND2_X1 U70 ( .A1(D[31]), .A2(n106), .ZN(n64) );
  BUF_X1 U71 ( .A(n73), .Z(n113) );
  BUF_X1 U72 ( .A(n73), .Z(n112) );
  BUF_X1 U73 ( .A(n73), .Z(n114) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n111) );
endmodule


module D_Reg_generic_N5_2 ( D, CLK, RESET, ENABLE, Q );
  input [4:0] D;
  output [4:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, net56157, net56158, net56159, net56160, net56161,
         n6, n7, n8, n9, n10, n12;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(CLK), .RN(RESET), .Q(Q[4]), .QN(net56161)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(CLK), .RN(RESET), .Q(Q[3]), .QN(net56160)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(CLK), .RN(RESET), .Q(Q[2]), .QN(net56159)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(CLK), .RN(RESET), .Q(Q[1]), .QN(net56158)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(CLK), .RN(RESET), .Q(Q[0]), .QN(net56157)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n12) );
  OAI21_X1 U3 ( .B1(net56158), .B2(n12), .A(n7), .ZN(n4) );
  NAND2_X1 U4 ( .A1(D[1]), .A2(n12), .ZN(n7) );
  OAI21_X1 U5 ( .B1(net56159), .B2(n12), .A(n8), .ZN(n3) );
  NAND2_X1 U6 ( .A1(D[2]), .A2(n12), .ZN(n8) );
  OAI21_X1 U7 ( .B1(net56160), .B2(n12), .A(n9), .ZN(n2) );
  NAND2_X1 U8 ( .A1(D[3]), .A2(n12), .ZN(n9) );
  OAI21_X1 U9 ( .B1(net56161), .B2(n12), .A(n10), .ZN(n1) );
  NAND2_X1 U10 ( .A1(D[4]), .A2(n12), .ZN(n10) );
  OAI21_X1 U11 ( .B1(net56157), .B2(n12), .A(n6), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n12), .A2(D[0]), .ZN(n6) );
endmodule


module D_Reg_generic_N32_3 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55837, net55838, net55839, net55840, net55841, net55842,
         net55843, net55844, net55845, net55846, net55847, net55848, net55849,
         net55850, net55851, net55852, net55853, net55854, net55855, net55856,
         net55857, net55858, net55859, net55860, net55861, net55862, net55863,
         net55864, net55865, net55866, net55867, net55868, n73, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n106, n107, n108, n109, n110, n111, n112, n113, n114;
  assign n73 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n114), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n112), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n114), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n112), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n114), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n112), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n112), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n112), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n114), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n112), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n112), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n112), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n114), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n113), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n113), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n113), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n112), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n113), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n113), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n113), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n113), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n113), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n114), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n112), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n114), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n112), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n113), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n112), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n113), .Q(Q[3]), .QN(net55840)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n113), .Q(Q[2]), .QN(net55839)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n113), .Q(Q[1]), .QN(net55838)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n114), .Q(Q[0]), .QN(net55837)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n106) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n108) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n110) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n109) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n107) );
  OAI21_X1 U7 ( .B1(net55860), .B2(n109), .A(n33), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n111), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U9 ( .B1(net55837), .B2(n109), .A(n39), .ZN(n32) );
  OAI21_X1 U10 ( .B1(net55857), .B2(n111), .A(n61), .ZN(n12) );
  NAND2_X1 U11 ( .A1(D[20]), .A2(n106), .ZN(n61) );
  OAI21_X1 U12 ( .B1(net55858), .B2(n111), .A(n62), .ZN(n11) );
  NAND2_X1 U13 ( .A1(D[21]), .A2(n106), .ZN(n62) );
  OAI21_X1 U14 ( .B1(net55859), .B2(n111), .A(n63), .ZN(n10) );
  NAND2_X1 U15 ( .A1(D[22]), .A2(n106), .ZN(n63) );
  OAI21_X1 U16 ( .B1(net55853), .B2(n110), .A(n57), .ZN(n16) );
  NAND2_X1 U17 ( .A1(D[16]), .A2(n106), .ZN(n57) );
  OAI21_X1 U18 ( .B1(net55854), .B2(n110), .A(n58), .ZN(n15) );
  NAND2_X1 U19 ( .A1(D[17]), .A2(n106), .ZN(n58) );
  OAI21_X1 U20 ( .B1(net55855), .B2(n110), .A(n59), .ZN(n14) );
  NAND2_X1 U21 ( .A1(D[18]), .A2(n106), .ZN(n59) );
  OAI21_X1 U22 ( .B1(net55856), .B2(n110), .A(n60), .ZN(n13) );
  NAND2_X1 U23 ( .A1(D[19]), .A2(n106), .ZN(n60) );
  OAI21_X1 U24 ( .B1(net55861), .B2(n108), .A(n34), .ZN(n8) );
  NAND2_X1 U25 ( .A1(D[24]), .A2(n106), .ZN(n34) );
  OAI21_X1 U26 ( .B1(net55862), .B2(n108), .A(n35), .ZN(n7) );
  NAND2_X1 U27 ( .A1(D[25]), .A2(n106), .ZN(n35) );
  OAI21_X1 U28 ( .B1(net55863), .B2(n109), .A(n36), .ZN(n6) );
  NAND2_X1 U29 ( .A1(D[26]), .A2(n106), .ZN(n36) );
  OAI21_X1 U30 ( .B1(net55864), .B2(n108), .A(n37), .ZN(n5) );
  NAND2_X1 U31 ( .A1(D[27]), .A2(n106), .ZN(n37) );
  OAI21_X1 U32 ( .B1(net55868), .B2(n109), .A(n64), .ZN(n1) );
  NAND2_X1 U33 ( .A1(D[31]), .A2(n106), .ZN(n64) );
  OAI21_X1 U34 ( .B1(net55841), .B2(n109), .A(n44), .ZN(n28) );
  NAND2_X1 U35 ( .A1(D[4]), .A2(n108), .ZN(n44) );
  OAI21_X1 U36 ( .B1(net55842), .B2(n109), .A(n45), .ZN(n27) );
  NAND2_X1 U37 ( .A1(D[5]), .A2(n108), .ZN(n45) );
  OAI21_X1 U38 ( .B1(net55843), .B2(n109), .A(n46), .ZN(n26) );
  NAND2_X1 U39 ( .A1(D[6]), .A2(n108), .ZN(n46) );
  OAI21_X1 U40 ( .B1(net55844), .B2(n109), .A(n47), .ZN(n25) );
  NAND2_X1 U41 ( .A1(D[7]), .A2(n108), .ZN(n47) );
  OAI21_X1 U42 ( .B1(net55845), .B2(n109), .A(n48), .ZN(n24) );
  NAND2_X1 U43 ( .A1(D[8]), .A2(n108), .ZN(n48) );
  OAI21_X1 U44 ( .B1(net55846), .B2(n110), .A(n49), .ZN(n23) );
  NAND2_X1 U45 ( .A1(D[9]), .A2(n108), .ZN(n49) );
  OAI21_X1 U46 ( .B1(net55866), .B2(n109), .A(n42), .ZN(n3) );
  NAND2_X1 U47 ( .A1(D[29]), .A2(n108), .ZN(n42) );
  OAI21_X1 U48 ( .B1(net55838), .B2(n108), .A(n40), .ZN(n31) );
  NAND2_X1 U49 ( .A1(D[1]), .A2(n107), .ZN(n40) );
  OAI21_X1 U50 ( .B1(net55839), .B2(n109), .A(n41), .ZN(n30) );
  NAND2_X1 U51 ( .A1(D[2]), .A2(n107), .ZN(n41) );
  OAI21_X1 U52 ( .B1(net55840), .B2(n109), .A(n43), .ZN(n29) );
  NAND2_X1 U53 ( .A1(D[3]), .A2(n107), .ZN(n43) );
  OAI21_X1 U54 ( .B1(net55847), .B2(n110), .A(n50), .ZN(n22) );
  NAND2_X1 U55 ( .A1(D[10]), .A2(n107), .ZN(n50) );
  OAI21_X1 U56 ( .B1(net55848), .B2(n110), .A(n51), .ZN(n21) );
  NAND2_X1 U57 ( .A1(D[11]), .A2(n107), .ZN(n51) );
  OAI21_X1 U58 ( .B1(net55849), .B2(n110), .A(n52), .ZN(n20) );
  NAND2_X1 U59 ( .A1(D[12]), .A2(n107), .ZN(n52) );
  OAI21_X1 U60 ( .B1(net55850), .B2(n110), .A(n54), .ZN(n19) );
  NAND2_X1 U61 ( .A1(D[13]), .A2(n107), .ZN(n54) );
  OAI21_X1 U62 ( .B1(net55851), .B2(n110), .A(n55), .ZN(n18) );
  NAND2_X1 U63 ( .A1(D[14]), .A2(n107), .ZN(n55) );
  OAI21_X1 U64 ( .B1(net55852), .B2(n110), .A(n56), .ZN(n17) );
  NAND2_X1 U65 ( .A1(D[15]), .A2(n107), .ZN(n56) );
  OAI21_X1 U66 ( .B1(net55865), .B2(n108), .A(n38), .ZN(n4) );
  NAND2_X1 U67 ( .A1(D[28]), .A2(n107), .ZN(n38) );
  OAI21_X1 U68 ( .B1(net55867), .B2(n110), .A(n53), .ZN(n2) );
  NAND2_X1 U69 ( .A1(D[30]), .A2(n107), .ZN(n53) );
  BUF_X1 U70 ( .A(n73), .Z(n113) );
  BUF_X1 U71 ( .A(n73), .Z(n112) );
  BUF_X1 U72 ( .A(n73), .Z(n114) );
  NAND2_X1 U73 ( .A1(D[0]), .A2(n107), .ZN(n39) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n111) );
endmodule


module D_Reg_generic_N32_4 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n49, net229340, net229338, net239847, net240147,
         net240375, net241423, net242614, net242616, net239809, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103;
  assign n49 = RESET;

  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n101), .Q(Q[26]) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n101), .Q(Q[25]) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n101), .Q(Q[24]) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n103), .Q(Q[23]) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n101), .Q(Q[22]) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n101), .Q(Q[21]) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n101), .Q(Q[20]) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n103), .Q(Q[19]) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n102), .Q(Q[18]) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n102), .Q(Q[17]) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n102), .Q(Q[16]) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n101), .Q(Q[15]) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n102), .Q(Q[14]) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n102), .Q(Q[13]) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n102), .Q(Q[12]) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n102), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n102), .Q(Q[10]) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n103), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n101), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n102), .Q(Q[5]) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n102), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n102), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n102), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n103), .Q(Q[0]) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n101), .Q(Q[4]) );
  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n103), .Q(Q[31]), .QN(n33) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n101), .Q(Q[28]) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n49), .Q(Q[8]) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n49), .Q(Q[9]) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n49), .Q(Q[27]) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n49), .Q(Q[30]) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n103), .Q(Q[29]) );
  NAND2_X2 U2 ( .A1(Q[30]), .A2(net242614), .ZN(n94) );
  BUF_X2 U3 ( .A(ENABLE), .Z(net229338) );
  NAND2_X1 U4 ( .A1(D[28]), .A2(ENABLE), .ZN(n99) );
  NAND2_X1 U5 ( .A1(D[31]), .A2(ENABLE), .ZN(n92) );
  NAND2_X1 U6 ( .A1(n92), .A2(net239809), .ZN(n1) );
  OR2_X1 U7 ( .A1(net229338), .A2(n33), .ZN(net239809) );
  BUF_X2 U8 ( .A(ENABLE), .Z(net229340) );
  NAND2_X1 U9 ( .A1(D[30]), .A2(net242616), .ZN(n93) );
  NAND2_X1 U10 ( .A1(n93), .A2(n94), .ZN(n2) );
  INV_X1 U11 ( .A(net242614), .ZN(net242616) );
  INV_X1 U12 ( .A(net229338), .ZN(net242614) );
  NAND2_X1 U13 ( .A1(D[29]), .A2(net241423), .ZN(n95) );
  NAND2_X2 U14 ( .A1(Q[29]), .A2(net239847), .ZN(n96) );
  NAND2_X1 U15 ( .A1(n95), .A2(n96), .ZN(n3) );
  INV_X1 U16 ( .A(net239847), .ZN(net241423) );
  INV_X1 U17 ( .A(net229338), .ZN(net239847) );
  NAND2_X1 U18 ( .A1(D[27]), .A2(net240375), .ZN(n97) );
  NAND2_X2 U19 ( .A1(Q[27]), .A2(net240147), .ZN(n98) );
  NAND2_X1 U20 ( .A1(n97), .A2(n98), .ZN(n5) );
  INV_X1 U21 ( .A(net240147), .ZN(net240375) );
  INV_X1 U22 ( .A(net229338), .ZN(net240147) );
  NAND2_X2 U23 ( .A1(Q[28]), .A2(net239847), .ZN(n100) );
  NAND2_X1 U24 ( .A1(n99), .A2(n100), .ZN(n4) );
  BUF_X1 U25 ( .A(n49), .Z(n102) );
  BUF_X1 U26 ( .A(n49), .Z(n101) );
  BUF_X1 U27 ( .A(n49), .Z(n103) );
  MUX2_X1 U28 ( .A(Q[4]), .B(D[4]), .S(net229338), .Z(n28) );
  MUX2_X1 U29 ( .A(Q[0]), .B(D[0]), .S(net229338), .Z(n32) );
  MUX2_X1 U30 ( .A(Q[1]), .B(D[1]), .S(net229338), .Z(n31) );
  MUX2_X1 U31 ( .A(Q[2]), .B(D[2]), .S(net229338), .Z(n30) );
  MUX2_X1 U32 ( .A(Q[3]), .B(D[3]), .S(net229338), .Z(n29) );
  MUX2_X1 U33 ( .A(Q[5]), .B(D[5]), .S(net229338), .Z(n27) );
  MUX2_X1 U34 ( .A(Q[6]), .B(D[6]), .S(net229338), .Z(n26) );
  MUX2_X1 U35 ( .A(Q[7]), .B(D[7]), .S(net229338), .Z(n25) );
  MUX2_X1 U36 ( .A(Q[8]), .B(D[8]), .S(net229338), .Z(n24) );
  MUX2_X1 U37 ( .A(Q[9]), .B(D[9]), .S(net229338), .Z(n23) );
  MUX2_X1 U38 ( .A(Q[10]), .B(D[10]), .S(net229338), .Z(n22) );
  MUX2_X1 U39 ( .A(Q[11]), .B(D[11]), .S(net229340), .Z(n21) );
  MUX2_X1 U40 ( .A(Q[12]), .B(D[12]), .S(net229340), .Z(n20) );
  MUX2_X1 U41 ( .A(Q[13]), .B(D[13]), .S(net229340), .Z(n19) );
  MUX2_X1 U42 ( .A(Q[14]), .B(D[14]), .S(net229340), .Z(n18) );
  MUX2_X1 U43 ( .A(Q[15]), .B(D[15]), .S(net229340), .Z(n17) );
  MUX2_X1 U44 ( .A(Q[16]), .B(D[16]), .S(net229340), .Z(n16) );
  MUX2_X1 U45 ( .A(Q[17]), .B(D[17]), .S(net229340), .Z(n15) );
  MUX2_X1 U46 ( .A(Q[18]), .B(D[18]), .S(net229340), .Z(n14) );
  MUX2_X1 U47 ( .A(Q[19]), .B(D[19]), .S(net229340), .Z(n13) );
  MUX2_X1 U48 ( .A(Q[20]), .B(D[20]), .S(net229340), .Z(n12) );
  MUX2_X1 U49 ( .A(Q[21]), .B(D[21]), .S(net229340), .Z(n11) );
  MUX2_X1 U50 ( .A(Q[22]), .B(D[22]), .S(net229340), .Z(n10) );
  MUX2_X1 U51 ( .A(Q[23]), .B(D[23]), .S(net229340), .Z(n9) );
  MUX2_X1 U52 ( .A(Q[24]), .B(D[24]), .S(net229340), .Z(n8) );
  MUX2_X1 U53 ( .A(Q[25]), .B(D[25]), .S(net229340), .Z(n7) );
  MUX2_X1 U54 ( .A(Q[26]), .B(D[26]), .S(net229340), .Z(n6) );
endmodule


module D_Reg_generic_N32_5 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55837, net55838, net55839, net55840, net55841, net55842,
         net55843, net55844, net55845, net55846, net55847, net55848, net55849,
         net55850, net55851, net55852, net55853, net55854, net55855, net55856,
         net55857, net55858, net55859, net55860, net55861, net55862, net55863,
         net55864, net55865, net55866, net55867, net55868, n73, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n106, n107, n108, n109, n110, n111, n112, n113, n114;
  assign n73 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n114), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n112), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n114), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n112), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n114), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n112), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n112), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n112), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n114), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n112), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n112), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n112), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n114), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n113), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n113), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n113), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n112), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n113), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n113), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n113), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n113), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n113), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n114), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n112), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n114), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n112), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n113), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n112), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n113), .Q(Q[3]), .QN(net55840)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n113), .Q(Q[2]), .QN(net55839)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n113), .Q(Q[1]), .QN(net55838)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n114), .Q(Q[0]), .QN(net55837)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n106) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n108) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n110) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n109) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n107) );
  OAI21_X1 U7 ( .B1(net55860), .B2(n109), .A(n33), .ZN(n9) );
  NAND2_X1 U8 ( .A1(n111), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U9 ( .B1(net55839), .B2(n109), .A(n41), .ZN(n30) );
  OAI21_X1 U10 ( .B1(net55857), .B2(n111), .A(n61), .ZN(n12) );
  NAND2_X1 U11 ( .A1(D[20]), .A2(n106), .ZN(n61) );
  OAI21_X1 U12 ( .B1(net55858), .B2(n111), .A(n62), .ZN(n11) );
  NAND2_X1 U13 ( .A1(D[21]), .A2(n106), .ZN(n62) );
  OAI21_X1 U14 ( .B1(net55859), .B2(n111), .A(n63), .ZN(n10) );
  NAND2_X1 U15 ( .A1(D[22]), .A2(n106), .ZN(n63) );
  OAI21_X1 U16 ( .B1(net55853), .B2(n110), .A(n57), .ZN(n16) );
  NAND2_X1 U17 ( .A1(D[16]), .A2(n106), .ZN(n57) );
  OAI21_X1 U18 ( .B1(net55854), .B2(n110), .A(n58), .ZN(n15) );
  NAND2_X1 U19 ( .A1(D[17]), .A2(n106), .ZN(n58) );
  OAI21_X1 U20 ( .B1(net55855), .B2(n110), .A(n59), .ZN(n14) );
  NAND2_X1 U21 ( .A1(D[18]), .A2(n106), .ZN(n59) );
  OAI21_X1 U22 ( .B1(net55856), .B2(n110), .A(n60), .ZN(n13) );
  NAND2_X1 U23 ( .A1(D[19]), .A2(n106), .ZN(n60) );
  OAI21_X1 U24 ( .B1(net55861), .B2(n108), .A(n34), .ZN(n8) );
  NAND2_X1 U25 ( .A1(D[24]), .A2(n106), .ZN(n34) );
  OAI21_X1 U26 ( .B1(net55862), .B2(n108), .A(n35), .ZN(n7) );
  NAND2_X1 U27 ( .A1(D[25]), .A2(n106), .ZN(n35) );
  OAI21_X1 U28 ( .B1(net55863), .B2(n109), .A(n36), .ZN(n6) );
  NAND2_X1 U29 ( .A1(D[26]), .A2(n106), .ZN(n36) );
  OAI21_X1 U30 ( .B1(net55864), .B2(n108), .A(n37), .ZN(n5) );
  NAND2_X1 U31 ( .A1(D[27]), .A2(n106), .ZN(n37) );
  OAI21_X1 U32 ( .B1(net55868), .B2(n109), .A(n64), .ZN(n1) );
  NAND2_X1 U33 ( .A1(D[31]), .A2(n106), .ZN(n64) );
  OAI21_X1 U34 ( .B1(net55841), .B2(n109), .A(n44), .ZN(n28) );
  NAND2_X1 U35 ( .A1(D[4]), .A2(n108), .ZN(n44) );
  OAI21_X1 U36 ( .B1(net55842), .B2(n109), .A(n45), .ZN(n27) );
  NAND2_X1 U37 ( .A1(D[5]), .A2(n108), .ZN(n45) );
  OAI21_X1 U38 ( .B1(net55843), .B2(n109), .A(n46), .ZN(n26) );
  NAND2_X1 U39 ( .A1(D[6]), .A2(n108), .ZN(n46) );
  OAI21_X1 U40 ( .B1(net55844), .B2(n109), .A(n47), .ZN(n25) );
  NAND2_X1 U41 ( .A1(D[7]), .A2(n108), .ZN(n47) );
  OAI21_X1 U42 ( .B1(net55845), .B2(n109), .A(n48), .ZN(n24) );
  NAND2_X1 U43 ( .A1(D[8]), .A2(n108), .ZN(n48) );
  OAI21_X1 U44 ( .B1(net55846), .B2(n110), .A(n49), .ZN(n23) );
  NAND2_X1 U45 ( .A1(D[9]), .A2(n108), .ZN(n49) );
  OAI21_X1 U46 ( .B1(net55866), .B2(n109), .A(n42), .ZN(n3) );
  NAND2_X1 U47 ( .A1(D[29]), .A2(n108), .ZN(n42) );
  OAI21_X1 U48 ( .B1(net55837), .B2(n109), .A(n39), .ZN(n32) );
  NAND2_X1 U49 ( .A1(D[0]), .A2(n107), .ZN(n39) );
  OAI21_X1 U50 ( .B1(net55838), .B2(n108), .A(n40), .ZN(n31) );
  NAND2_X1 U51 ( .A1(D[1]), .A2(n107), .ZN(n40) );
  OAI21_X1 U52 ( .B1(net55840), .B2(n109), .A(n43), .ZN(n29) );
  NAND2_X1 U53 ( .A1(D[3]), .A2(n107), .ZN(n43) );
  OAI21_X1 U54 ( .B1(net55847), .B2(n110), .A(n50), .ZN(n22) );
  NAND2_X1 U55 ( .A1(D[10]), .A2(n107), .ZN(n50) );
  OAI21_X1 U56 ( .B1(net55848), .B2(n110), .A(n51), .ZN(n21) );
  NAND2_X1 U57 ( .A1(D[11]), .A2(n107), .ZN(n51) );
  OAI21_X1 U58 ( .B1(net55849), .B2(n110), .A(n52), .ZN(n20) );
  NAND2_X1 U59 ( .A1(D[12]), .A2(n107), .ZN(n52) );
  OAI21_X1 U60 ( .B1(net55850), .B2(n110), .A(n54), .ZN(n19) );
  NAND2_X1 U61 ( .A1(D[13]), .A2(n107), .ZN(n54) );
  OAI21_X1 U62 ( .B1(net55851), .B2(n110), .A(n55), .ZN(n18) );
  NAND2_X1 U63 ( .A1(D[14]), .A2(n107), .ZN(n55) );
  OAI21_X1 U64 ( .B1(net55852), .B2(n110), .A(n56), .ZN(n17) );
  NAND2_X1 U65 ( .A1(D[15]), .A2(n107), .ZN(n56) );
  OAI21_X1 U66 ( .B1(net55865), .B2(n108), .A(n38), .ZN(n4) );
  NAND2_X1 U67 ( .A1(D[28]), .A2(n107), .ZN(n38) );
  OAI21_X1 U68 ( .B1(net55867), .B2(n110), .A(n53), .ZN(n2) );
  NAND2_X1 U69 ( .A1(D[30]), .A2(n107), .ZN(n53) );
  BUF_X1 U70 ( .A(n73), .Z(n113) );
  BUF_X1 U71 ( .A(n73), .Z(n112) );
  BUF_X1 U72 ( .A(n73), .Z(n114) );
  NAND2_X1 U73 ( .A1(D[2]), .A2(n107), .ZN(n41) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n111) );
endmodule


module ALU_N32 ( FUNC, Sign, AddrComp, DATA1, DATA2, OUTALU );
  input [4:0] FUNC;
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  input Sign, AddrComp;
  wire   Sub, L_A, L_R, S_R, Cout, Sign_OF, Unsign_OF, AneB, AeqB, AgtB, AgeB,
         AltB, AleB, \Comp_ext[0] , OvFl, \Over[31] , n50, n53, n55, n58, n59,
         n63, n65, n69, n70, n75, n77, n78, n79, n80, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236;
  wire   [2:0] Comp_Sel;
  wire   [2:0] Out_Sel;
  wire   [31:0] And_Out;
  wire   [31:0] Or_Out;
  wire   [31:0] Xor_Out;
  wire   [31:0] Add_Out;
  wire   [31:0] Shift_Out;
  wire   [31:0] Mul_Out;
  wire   [31:0] Add_Ok;
  assign n50 = DATA1[4];
  assign n53 = DATA1[8];
  assign n55 = DATA1[6];
  assign n58 = DATA1[3];
  assign n59 = DATA2[3];
  assign n63 = DATA1[7];
  assign n65 = DATA1[0];
  assign n69 = DATA1[5];
  assign n70 = DATA1[2];
  assign n75 = DATA1[9];
  assign n77 = DATA2[0];
  assign n78 = DATA1[1];
  assign n79 = DATA2[2];
  assign n80 = DATA2[1];
  assign n87 = DATA1[15];
  assign n88 = DATA1[10];
  assign n89 = DATA1[11];
  assign n90 = DATA1[12];
  assign n91 = DATA1[13];
  assign n92 = DATA1[16];
  assign n93 = DATA1[20];
  assign n94 = DATA1[21];
  assign n95 = DATA1[22];
  assign n96 = DATA1[23];
  assign n97 = DATA1[24];
  assign n98 = DATA1[25];
  assign n99 = DATA1[26];

  and_gen_N32 AND_OP ( .A({DATA1[31:27], n198, n197, n196, n96, n195, n94, 
        n194, DATA1[19:17], n92, n189, DATA1[14], n193, n192, n191, n88, n75, 
        n152, n164, n148, n158, n162, n181, n166, n182, n169}), .B({
        DATA2[31:5], n150, n159, n184, n175, n172}), .C(And_Out) );
  or_gen_N32 OR_OP ( .A({DATA1[31:27], n198, n197, n196, n96, n195, n94, n194, 
        DATA1[19:17], n92, n189, DATA1[14], n193, n192, n191, n88, n75, n152, 
        n165, n55, n158, n161, n190, n166, n183, n169}), .B({DATA2[31:5], n150, 
        n159, n184, n175, n172}), .C(Or_Out) );
  xor_gen_N32_0 XOR_OP ( .A({DATA1[31:27], n198, n197, n196, n96, n195, n94, 
        n194, DATA1[19:17], n92, n189, DATA1[14], n193, n192, n191, n88, n75, 
        n152, n164, n55, n158, n161, n181, n166, n182, n169}), .B({DATA2[31:5], 
        n150, n159, n184, n175, n172}), .C(Xor_Out) );
  Add_gen_N32 ADDER ( .A({DATA1[31:27], n198, n197, n196, n96, n195, n94, n194, 
        DATA1[19:17], n92, n189, DATA1[14], n193, n192, n191, n88, n75, n152, 
        n164, n55, n69, n154, n181, n166, n183, n168}), .B({DATA2[31:5], n150, 
        n59, n184, n175, n172}), .sub(Sub), .S(Add_Out), .Co(Cout), .Sign_OF(
        Sign_OF), .Unsign_OF(Unsign_OF) );
  SHIFTER_GENERIC_N32 SH_ROT ( .A({DATA1[31:27], n198, n197, n196, n96, n195, 
        n94, n194, DATA1[19:17], n92, n189, DATA1[14], n193, n192, n191, n88, 
        n75, n152, n165, n55, n156, n154, n190, n166, n173, n168}), .B({n150, 
        n59, n170, n175, n172}), .LOGIC_ARITH(L_A), .LEFT_RIGHT(L_R), 
        .SHIFT_ROTATE(S_R), .OUTPUT(Shift_Out) );
  Comparator_Nbit32 COMP ( .Diff(Add_Out), .Cout(Cout), .Sign(Sign), .a(
        DATA1[31]), .b(DATA2[31]), .Ne(AneB), .Eq(AeqB), .Gt(AgtB), .Ge(AgeB), 
        .Lt(AltB), .Le(AleB) );
  Boothmul_N16 MUL ( .A({n189, DATA1[14], n193, n192, n191, n88, n75, n53, 
        n188, n55, n69, n50, n190, n70, n78, n65}), .B({DATA2[15:4], n59, n79, 
        n80, n77}), .P(Mul_Out) );
  mux81_logic MuxComp ( .A(AneB), .B(AeqB), .C(AgtB), .D(AgeB), .E(AltB), .F(
        AleB), .G(1'b0), .H(1'b0), .S(Comp_Sel), .Y(\Comp_ext[0] ) );
  MUX21_919 OF_Detect ( .A(Unsign_OF), .B(Sign_OF), .S(Sign), .Y(OvFl) );
  MUX21_GENERIC_N32_11 OF_Manage ( .A(Add_Out), .B({\Over[31] , n185, n185, 
        n185, n185, n185, n186, n185, n185, n185, n185, n185, n185, n186, n186, 
        n186, n186, n186, n186, n186, n186, n186, n186, n186, n186, n187, n187, 
        n187, n187, n187, n187, n185}), .S(n179), .Y(Add_Ok) );
  mux81_generic_N32 MuxOut ( .A(And_Out), .B(Or_Out), .C(Xor_Out), .D(Add_Ok), 
        .E(Shift_Out), .F({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \Comp_ext[0] }), .G(Mul_Out), .H({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .S(Out_Sel), .Y(OUTALU) );
  CLKBUF_X1 U2 ( .A(n55), .Z(n148) );
  BUF_X4 U3 ( .A(n58), .Z(n190) );
  INV_X8 U4 ( .A(n171), .ZN(n172) );
  CLKBUF_X1 U5 ( .A(n70), .Z(n166) );
  INV_X1 U6 ( .A(DATA2[4]), .ZN(n149) );
  INV_X2 U7 ( .A(n149), .ZN(n150) );
  BUF_X4 U8 ( .A(n89), .Z(n191) );
  BUF_X4 U9 ( .A(n90), .Z(n192) );
  INV_X1 U10 ( .A(n53), .ZN(n151) );
  INV_X2 U11 ( .A(n151), .ZN(n152) );
  INV_X1 U12 ( .A(n50), .ZN(n153) );
  INV_X2 U13 ( .A(n153), .ZN(n154) );
  INV_X1 U14 ( .A(n69), .ZN(n155) );
  INV_X2 U15 ( .A(n155), .ZN(n156) );
  CLKBUF_X1 U16 ( .A(n78), .Z(n157) );
  CLKBUF_X1 U17 ( .A(n156), .Z(n158) );
  CLKBUF_X1 U18 ( .A(n59), .Z(n159) );
  CLKBUF_X1 U19 ( .A(n80), .Z(n160) );
  CLKBUF_X1 U20 ( .A(n154), .Z(n161) );
  CLKBUF_X1 U21 ( .A(n154), .Z(n162) );
  CLKBUF_X1 U22 ( .A(n157), .Z(n163) );
  BUF_X4 U23 ( .A(n91), .Z(n193) );
  CLKBUF_X1 U24 ( .A(n63), .Z(n165) );
  CLKBUF_X1 U25 ( .A(n63), .Z(n164) );
  CLKBUF_X1 U26 ( .A(n79), .Z(n170) );
  INV_X1 U27 ( .A(n65), .ZN(n167) );
  INV_X2 U28 ( .A(n167), .ZN(n168) );
  BUF_X4 U29 ( .A(n87), .Z(n189) );
  CLKBUF_X1 U30 ( .A(n168), .Z(n169) );
  INV_X1 U31 ( .A(n77), .ZN(n171) );
  CLKBUF_X1 U32 ( .A(n163), .Z(n173) );
  INV_X1 U33 ( .A(n160), .ZN(n174) );
  INV_X4 U34 ( .A(n174), .ZN(n175) );
  BUF_X1 U35 ( .A(n98), .Z(n197) );
  BUF_X1 U36 ( .A(n99), .Z(n198) );
  BUF_X1 U37 ( .A(n97), .Z(n196) );
  BUF_X1 U38 ( .A(n93), .Z(n194) );
  BUF_X1 U39 ( .A(n95), .Z(n195) );
  NAND2_X1 U40 ( .A1(n178), .A2(n218), .ZN(n232) );
  INV_X1 U41 ( .A(Sub), .ZN(n185) );
  INV_X1 U42 ( .A(Sub), .ZN(n186) );
  NAND2_X1 U43 ( .A1(n204), .A2(n217), .ZN(Sub) );
  NAND2_X1 U44 ( .A1(n208), .A2(n220), .ZN(n221) );
  AND2_X1 U45 ( .A1(n236), .A2(n199), .ZN(n176) );
  NAND2_X1 U46 ( .A1(n200), .A2(n176), .ZN(n220) );
  NOR2_X1 U47 ( .A1(n232), .A2(n231), .ZN(n235) );
  NOR2_X1 U48 ( .A1(n232), .A2(n223), .ZN(n222) );
  OAI21_X1 U49 ( .B1(n205), .B2(n230), .A(n177), .ZN(n216) );
  AND2_X1 U50 ( .A1(n211), .A2(n206), .ZN(n177) );
  NAND2_X1 U51 ( .A1(n211), .A2(n221), .ZN(n218) );
  AND3_X1 U52 ( .A1(n217), .A2(n216), .A3(n227), .ZN(n178) );
  NOR2_X1 U53 ( .A1(n231), .A2(n223), .ZN(n224) );
  AND2_X1 U54 ( .A1(OvFl), .A2(n229), .ZN(n179) );
  NAND2_X1 U55 ( .A1(n202), .A2(n201), .ZN(n223) );
  NAND2_X1 U56 ( .A1(n210), .A2(n219), .ZN(n231) );
  AND2_X1 U57 ( .A1(FUNC[3]), .A2(FUNC[2]), .ZN(n180) );
  NAND2_X1 U58 ( .A1(n200), .A2(FUNC[1]), .ZN(n207) );
  CLKBUF_X1 U59 ( .A(n157), .Z(n183) );
  CLKBUF_X1 U60 ( .A(n163), .Z(n182) );
  CLKBUF_X1 U61 ( .A(n58), .Z(n181) );
  CLKBUF_X1 U62 ( .A(n170), .Z(n184) );
  BUF_X4 U63 ( .A(n63), .Z(n188) );
  INV_X1 U64 ( .A(Sub), .ZN(n187) );
  INV_X1 U65 ( .A(FUNC[1]), .ZN(n199) );
  INV_X1 U66 ( .A(FUNC[4]), .ZN(n200) );
  NAND3_X1 U67 ( .A1(FUNC[0]), .A2(n199), .A3(n200), .ZN(n208) );
  INV_X1 U68 ( .A(FUNC[0]), .ZN(n236) );
  NAND2_X1 U69 ( .A1(n180), .A2(n221), .ZN(n202) );
  INV_X1 U70 ( .A(n207), .ZN(n230) );
  NAND2_X1 U71 ( .A1(FUNC[3]), .A2(n230), .ZN(n201) );
  INV_X1 U72 ( .A(n223), .ZN(n204) );
  INV_X1 U73 ( .A(n220), .ZN(n203) );
  INV_X1 U74 ( .A(FUNC[3]), .ZN(n211) );
  NAND3_X1 U75 ( .A1(FUNC[2]), .A2(n203), .A3(n211), .ZN(n217) );
  NAND2_X1 U76 ( .A1(FUNC[4]), .A2(n176), .ZN(n225) );
  INV_X1 U77 ( .A(n225), .ZN(n205) );
  INV_X1 U78 ( .A(FUNC[2]), .ZN(n206) );
  NAND3_X1 U79 ( .A1(FUNC[3]), .A2(n221), .A3(n206), .ZN(n210) );
  NAND2_X1 U80 ( .A1(n208), .A2(n207), .ZN(n209) );
  NAND3_X1 U81 ( .A1(FUNC[2]), .A2(n209), .A3(n211), .ZN(n219) );
  INV_X1 U82 ( .A(n231), .ZN(n215) );
  INV_X1 U83 ( .A(n218), .ZN(n213) );
  INV_X1 U84 ( .A(n216), .ZN(n212) );
  NOR2_X1 U85 ( .A1(n213), .A2(n212), .ZN(n214) );
  NAND3_X1 U86 ( .A1(n187), .A2(n215), .A3(n214), .ZN(n227) );
  INV_X1 U87 ( .A(n178), .ZN(Out_Sel[1]) );
  NAND2_X1 U88 ( .A1(n219), .A2(n222), .ZN(S_R) );
  NAND2_X1 U89 ( .A1(n220), .A2(n222), .ZN(L_R) );
  INV_X1 U90 ( .A(n221), .ZN(n234) );
  NAND3_X1 U91 ( .A1(FUNC[0]), .A2(n222), .A3(n234), .ZN(L_A) );
  NAND3_X1 U92 ( .A1(n225), .A2(n227), .A3(n224), .ZN(Out_Sel[2]) );
  NAND2_X1 U93 ( .A1(FUNC[0]), .A2(n177), .ZN(n226) );
  NAND3_X1 U94 ( .A1(n187), .A2(n227), .A3(n226), .ZN(Out_Sel[0]) );
  INV_X1 U95 ( .A(Sign), .ZN(n228) );
  XNOR2_X1 U96 ( .A(n185), .B(n228), .ZN(\Over[31] ) );
  INV_X1 U97 ( .A(AddrComp), .ZN(n229) );
  NAND2_X1 U98 ( .A1(n180), .A2(n230), .ZN(n233) );
  NAND2_X1 U99 ( .A1(n233), .A2(n235), .ZN(Comp_Sel[2]) );
  NAND2_X1 U100 ( .A1(n234), .A2(n235), .ZN(Comp_Sel[1]) );
  NAND2_X1 U101 ( .A1(n236), .A2(n235), .ZN(Comp_Sel[0]) );
endmodule


module mux41_generic_N32_2 ( A, B, C, D, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Y;

  wire   [31:0] ABto2;
  wire   [31:0] CDto2;

  MUX21_GENERIC_N32_14 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_GENERIC_N32_13 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_GENERIC_N32_12 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(Y) );
endmodule


module mux41_generic_N32_3 ( A, B, C, D, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Y;

  wire   [31:0] ABto2;
  wire   [31:0] CDto2;

  MUX21_GENERIC_N32_17 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_GENERIC_N32_16 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_GENERIC_N32_15 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(Y) );
endmodule


module Br_Comp_Nbit32 ( A, Br_cond, Taken );
  input [31:0] A;
  input [1:0] Br_cond;
  output Taken;
  wire   n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;

  XOR2_X1 U1 ( .A(n60), .B(Br_cond[0]), .Z(n62) );
  NOR2_X1 U2 ( .A1(A[23]), .A2(A[22]), .ZN(n41) );
  NOR2_X1 U3 ( .A1(A[21]), .A2(A[20]), .ZN(n40) );
  NOR2_X1 U4 ( .A1(A[19]), .A2(A[18]), .ZN(n39) );
  NOR2_X1 U5 ( .A1(A[17]), .A2(A[16]), .ZN(n38) );
  NAND4_X1 U6 ( .A1(n41), .A2(n40), .A3(n39), .A4(n38), .ZN(n47) );
  NOR2_X1 U7 ( .A1(A[31]), .A2(A[30]), .ZN(n45) );
  NOR2_X1 U8 ( .A1(A[29]), .A2(A[28]), .ZN(n44) );
  NOR2_X1 U9 ( .A1(A[27]), .A2(A[26]), .ZN(n43) );
  NOR2_X1 U10 ( .A1(A[25]), .A2(A[24]), .ZN(n42) );
  NAND4_X1 U11 ( .A1(n45), .A2(n44), .A3(n43), .A4(n42), .ZN(n46) );
  NOR2_X1 U12 ( .A1(n47), .A2(n46), .ZN(n59) );
  NOR2_X1 U13 ( .A1(A[7]), .A2(A[6]), .ZN(n51) );
  NOR2_X1 U14 ( .A1(A[5]), .A2(A[4]), .ZN(n50) );
  NOR2_X1 U15 ( .A1(A[3]), .A2(A[2]), .ZN(n49) );
  NOR2_X1 U16 ( .A1(A[1]), .A2(A[0]), .ZN(n48) );
  NAND4_X1 U17 ( .A1(n51), .A2(n50), .A3(n49), .A4(n48), .ZN(n57) );
  NOR2_X1 U18 ( .A1(A[15]), .A2(A[14]), .ZN(n55) );
  NOR2_X1 U19 ( .A1(A[13]), .A2(A[12]), .ZN(n54) );
  NOR2_X1 U20 ( .A1(A[11]), .A2(A[10]), .ZN(n53) );
  NOR2_X1 U21 ( .A1(A[9]), .A2(A[8]), .ZN(n52) );
  NAND4_X1 U22 ( .A1(n55), .A2(n54), .A3(n53), .A4(n52), .ZN(n56) );
  NOR2_X1 U23 ( .A1(n57), .A2(n56), .ZN(n58) );
  NAND2_X1 U24 ( .A1(n59), .A2(n58), .ZN(n60) );
  INV_X1 U25 ( .A(Br_cond[1]), .ZN(n61) );
  NOR2_X1 U26 ( .A1(n62), .A2(n61), .ZN(Taken) );
endmodule


module D_Reg_generic_N5_0 ( D, CLK, RESET, ENABLE, Q );
  input [4:0] D;
  output [4:0] Q;
  input CLK, RESET, ENABLE;
  wire   n11, n12, n13, n14, n15;

  DFFR_X1 \Q_reg[4]  ( .D(n15), .CK(CLK), .RN(RESET), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(n14), .CK(CLK), .RN(RESET), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(n13), .CK(CLK), .RN(RESET), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(n12), .CK(CLK), .RN(RESET), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(n11), .CK(CLK), .RN(RESET), .Q(Q[0]) );
  MUX2_X1 U2 ( .A(Q[0]), .B(D[0]), .S(ENABLE), .Z(n11) );
  MUX2_X1 U3 ( .A(Q[1]), .B(D[1]), .S(ENABLE), .Z(n12) );
  MUX2_X1 U4 ( .A(Q[2]), .B(D[2]), .S(ENABLE), .Z(n13) );
  MUX2_X1 U5 ( .A(Q[3]), .B(D[3]), .S(ENABLE), .Z(n14) );
  MUX2_X1 U6 ( .A(Q[4]), .B(D[4]), .S(ENABLE), .Z(n15) );
endmodule


module D_Reg_generic_N32_7 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55839, net55841, net55842, net55843, net55844, net55845,
         net55846, net55847, net55848, net55849, net55850, net55851, net55852,
         net55853, net55854, net55855, net55856, net55857, net55858, net55859,
         net55860, net55861, net55862, net55863, net55864, net55865, net55866,
         net55867, net55868, n124, n47, n81, n83, n84, n86, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123;
  assign n47 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n91), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n92), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n91), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n92), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n91), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n92), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n92), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n92), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n91), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n93), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n93), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n93), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n91), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n92), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n92), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n92), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n93), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n92), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n92), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n92), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n91), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n91), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n91), .Q(Q[9]), .QN(net55846) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n93), .Q(Q[8]), .QN(net55845) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n91), .Q(Q[7]), .QN(net55844) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n93), .Q(Q[6]), .QN(net55843) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n91), .Q(Q[5]), .QN(net55842) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n92), .Q(Q[4]), .QN(net55841) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n91), .Q(n124), .QN(n81) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n91), .Q(n83), .QN(net55839) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n47), .Q(n95), .QN(n84) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n47), .Q(n94), .QN(n86) );
  INV_X1 U2 ( .A(n81), .ZN(Q[3]) );
  INV_X1 U3 ( .A(n84), .ZN(Q[1]) );
  INV_X1 U4 ( .A(n86), .ZN(Q[0]) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n88) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n89) );
  BUF_X1 U7 ( .A(ENABLE), .Z(n90) );
  BUF_X1 U8 ( .A(n47), .Z(n92) );
  BUF_X1 U9 ( .A(n47), .Z(n91) );
  BUF_X1 U10 ( .A(n47), .Z(n93) );
  INV_X1 U11 ( .A(net55839), .ZN(Q[2]) );
  MUX2_X1 U12 ( .A(n94), .B(D[0]), .S(n88), .Z(n32) );
  MUX2_X1 U13 ( .A(n95), .B(D[1]), .S(n88), .Z(n31) );
  MUX2_X1 U14 ( .A(n83), .B(D[2]), .S(n88), .Z(n30) );
  MUX2_X1 U15 ( .A(n124), .B(D[3]), .S(n88), .Z(n29) );
  INV_X1 U16 ( .A(net55841), .ZN(n96) );
  MUX2_X1 U17 ( .A(n96), .B(D[4]), .S(n88), .Z(n28) );
  INV_X1 U18 ( .A(net55842), .ZN(n97) );
  MUX2_X1 U19 ( .A(n97), .B(D[5]), .S(n88), .Z(n27) );
  INV_X1 U20 ( .A(net55843), .ZN(n98) );
  MUX2_X1 U21 ( .A(n98), .B(D[6]), .S(n88), .Z(n26) );
  INV_X1 U22 ( .A(net55844), .ZN(n99) );
  MUX2_X1 U23 ( .A(n99), .B(D[7]), .S(n88), .Z(n25) );
  INV_X1 U24 ( .A(net55845), .ZN(n100) );
  MUX2_X1 U25 ( .A(n100), .B(D[8]), .S(n88), .Z(n24) );
  INV_X1 U26 ( .A(net55846), .ZN(n101) );
  MUX2_X1 U27 ( .A(n101), .B(D[9]), .S(n88), .Z(n23) );
  INV_X1 U28 ( .A(net55847), .ZN(n102) );
  MUX2_X1 U29 ( .A(n102), .B(D[10]), .S(n88), .Z(n22) );
  INV_X1 U30 ( .A(net55848), .ZN(n103) );
  MUX2_X1 U31 ( .A(n103), .B(D[11]), .S(n88), .Z(n21) );
  INV_X1 U32 ( .A(net55849), .ZN(n104) );
  MUX2_X1 U33 ( .A(n104), .B(D[12]), .S(n89), .Z(n20) );
  INV_X1 U34 ( .A(net55850), .ZN(n105) );
  MUX2_X1 U35 ( .A(n105), .B(D[13]), .S(n89), .Z(n19) );
  INV_X1 U36 ( .A(net55851), .ZN(n106) );
  MUX2_X1 U37 ( .A(n106), .B(D[14]), .S(n89), .Z(n18) );
  INV_X1 U38 ( .A(net55852), .ZN(n107) );
  MUX2_X1 U39 ( .A(n107), .B(D[15]), .S(n89), .Z(n17) );
  INV_X1 U40 ( .A(net55853), .ZN(n108) );
  MUX2_X1 U41 ( .A(n108), .B(D[16]), .S(n89), .Z(n16) );
  INV_X1 U42 ( .A(net55854), .ZN(n109) );
  MUX2_X1 U43 ( .A(n109), .B(D[17]), .S(n89), .Z(n15) );
  INV_X1 U44 ( .A(net55855), .ZN(n110) );
  MUX2_X1 U45 ( .A(n110), .B(D[18]), .S(n89), .Z(n14) );
  INV_X1 U46 ( .A(net55856), .ZN(n111) );
  MUX2_X1 U47 ( .A(n111), .B(D[19]), .S(n89), .Z(n13) );
  INV_X1 U48 ( .A(net55857), .ZN(n112) );
  MUX2_X1 U49 ( .A(n112), .B(D[20]), .S(n89), .Z(n12) );
  INV_X1 U50 ( .A(net55858), .ZN(n113) );
  MUX2_X1 U51 ( .A(n113), .B(D[21]), .S(n89), .Z(n11) );
  INV_X1 U52 ( .A(net55859), .ZN(n114) );
  MUX2_X1 U53 ( .A(n114), .B(D[22]), .S(n89), .Z(n10) );
  INV_X1 U54 ( .A(net55860), .ZN(n115) );
  MUX2_X1 U55 ( .A(n115), .B(D[23]), .S(n89), .Z(n9) );
  INV_X1 U56 ( .A(net55861), .ZN(n116) );
  MUX2_X1 U57 ( .A(n116), .B(D[24]), .S(n90), .Z(n8) );
  INV_X1 U58 ( .A(net55862), .ZN(n117) );
  MUX2_X1 U59 ( .A(n117), .B(D[25]), .S(n90), .Z(n7) );
  INV_X1 U60 ( .A(net55863), .ZN(n118) );
  MUX2_X1 U61 ( .A(n118), .B(D[26]), .S(n90), .Z(n6) );
  INV_X1 U62 ( .A(net55864), .ZN(n119) );
  MUX2_X1 U63 ( .A(n119), .B(D[27]), .S(n90), .Z(n5) );
  INV_X1 U64 ( .A(net55865), .ZN(n120) );
  MUX2_X1 U65 ( .A(n120), .B(D[28]), .S(n90), .Z(n4) );
  INV_X1 U66 ( .A(net55866), .ZN(n121) );
  MUX2_X1 U67 ( .A(n121), .B(D[29]), .S(n90), .Z(n3) );
  INV_X1 U68 ( .A(net55867), .ZN(n122) );
  MUX2_X1 U69 ( .A(n122), .B(D[30]), .S(n90), .Z(n2) );
  INV_X1 U70 ( .A(net55868), .ZN(n123) );
  MUX2_X1 U71 ( .A(n123), .B(D[31]), .S(n90), .Z(n1) );
endmodule


module D_Reg_generic_N32_8 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55840, net55841, net55842, net55843, net55844, net55845,
         net55846, net55847, net55848, net55849, net55850, net55851, net55852,
         net55853, net55854, net55855, net55856, net55857, net55858, net55859,
         net55860, net55861, net55862, net55863, net55864, net55865, net55866,
         net55867, net55868, n139, n85, n33, n34, n35, n36, n37, n38, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n118, n119, n127, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138;
  assign n85 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n136), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n138), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n136), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n138), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n136), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n138), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n137), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n137), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n136), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n137), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n137), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n137), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n136), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n137), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n137), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n136), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n138), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n136), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n137), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n137), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n136), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n136), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n136), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n138), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n136), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n137), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n137), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n137), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n85), .Q(n139), .QN(n127) );
  SDFFR_X1 \Q_reg[2]  ( .D(1'b0), .SI(n30), .SE(1'b1), .CK(CLK), .RN(n85), .Q(
        Q[2]) );
  SDFFR_X1 \Q_reg[1]  ( .D(1'b0), .SI(n31), .SE(1'b1), .CK(CLK), .RN(n85), .Q(
        Q[1]), .QN(n118) );
  SDFFR_X1 \Q_reg[3]  ( .D(1'b0), .SI(n29), .SE(1'b1), .CK(CLK), .RN(n136), 
        .Q(Q[3]), .QN(net55840) );
  INV_X1 U2 ( .A(n118), .ZN(n119) );
  INV_X1 U9 ( .A(n127), .ZN(Q[0]) );
  BUF_X1 U10 ( .A(n129), .Z(n131) );
  BUF_X1 U11 ( .A(n129), .Z(n132) );
  CLKBUF_X1 U12 ( .A(n129), .Z(n133) );
  BUF_X1 U13 ( .A(n130), .Z(n134) );
  BUF_X1 U14 ( .A(n130), .Z(n135) );
  BUF_X1 U15 ( .A(ENABLE), .Z(n129) );
  OAI21_X1 U16 ( .B1(net55860), .B2(n134), .A(n33), .ZN(n9) );
  NAND2_X1 U17 ( .A1(n135), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U18 ( .B1(net55840), .B2(n133), .A(n43), .ZN(n29) );
  NAND2_X1 U19 ( .A1(D[3]), .A2(n132), .ZN(n43) );
  OAI21_X1 U20 ( .B1(net55841), .B2(n133), .A(n44), .ZN(n28) );
  NAND2_X1 U21 ( .A1(D[4]), .A2(n132), .ZN(n44) );
  OAI21_X1 U22 ( .B1(net55861), .B2(n133), .A(n34), .ZN(n8) );
  NAND2_X1 U23 ( .A1(D[24]), .A2(n131), .ZN(n34) );
  OAI21_X1 U24 ( .B1(net55862), .B2(n133), .A(n35), .ZN(n7) );
  NAND2_X1 U25 ( .A1(D[25]), .A2(n131), .ZN(n35) );
  OAI21_X1 U26 ( .B1(net55863), .B2(n133), .A(n36), .ZN(n6) );
  NAND2_X1 U27 ( .A1(D[26]), .A2(n131), .ZN(n36) );
  OAI21_X1 U28 ( .B1(net55864), .B2(n133), .A(n37), .ZN(n5) );
  NAND2_X1 U29 ( .A1(D[27]), .A2(n131), .ZN(n37) );
  OAI21_X1 U30 ( .B1(net55865), .B2(n133), .A(n38), .ZN(n4) );
  NAND2_X1 U31 ( .A1(D[28]), .A2(n131), .ZN(n38) );
  OAI21_X1 U32 ( .B1(net55866), .B2(n133), .A(n42), .ZN(n3) );
  NAND2_X1 U33 ( .A1(D[29]), .A2(n132), .ZN(n42) );
  OAI21_X1 U34 ( .B1(net55844), .B2(n134), .A(n47), .ZN(n25) );
  NAND2_X1 U35 ( .A1(D[7]), .A2(n132), .ZN(n47) );
  OAI21_X1 U36 ( .B1(net55847), .B2(n134), .A(n50), .ZN(n22) );
  NAND2_X1 U37 ( .A1(D[10]), .A2(n132), .ZN(n50) );
  OAI21_X1 U38 ( .B1(net55848), .B2(n134), .A(n51), .ZN(n21) );
  NAND2_X1 U39 ( .A1(D[11]), .A2(n132), .ZN(n51) );
  OAI21_X1 U40 ( .B1(net55849), .B2(n134), .A(n52), .ZN(n20) );
  NAND2_X1 U41 ( .A1(D[12]), .A2(n132), .ZN(n52) );
  OAI21_X1 U42 ( .B1(net55850), .B2(n134), .A(n54), .ZN(n19) );
  NAND2_X1 U43 ( .A1(D[13]), .A2(n131), .ZN(n54) );
  OAI21_X1 U44 ( .B1(net55851), .B2(n134), .A(n55), .ZN(n18) );
  NAND2_X1 U45 ( .A1(D[14]), .A2(n132), .ZN(n55) );
  OAI21_X1 U46 ( .B1(net55867), .B2(n134), .A(n53), .ZN(n2) );
  NAND2_X1 U47 ( .A1(D[30]), .A2(n132), .ZN(n53) );
  OAI21_X1 U48 ( .B1(net55852), .B2(n135), .A(n56), .ZN(n17) );
  NAND2_X1 U49 ( .A1(D[15]), .A2(n132), .ZN(n56) );
  OAI21_X1 U50 ( .B1(net55853), .B2(n135), .A(n57), .ZN(n16) );
  NAND2_X1 U51 ( .A1(D[16]), .A2(n132), .ZN(n57) );
  OAI21_X1 U52 ( .B1(net55854), .B2(n135), .A(n58), .ZN(n15) );
  NAND2_X1 U53 ( .A1(D[17]), .A2(n132), .ZN(n58) );
  OAI21_X1 U54 ( .B1(net55855), .B2(n135), .A(n59), .ZN(n14) );
  NAND2_X1 U55 ( .A1(D[18]), .A2(n131), .ZN(n59) );
  OAI21_X1 U56 ( .B1(net55856), .B2(n135), .A(n60), .ZN(n13) );
  NAND2_X1 U57 ( .A1(D[19]), .A2(n131), .ZN(n60) );
  OAI21_X1 U58 ( .B1(net55857), .B2(n135), .A(n61), .ZN(n12) );
  NAND2_X1 U59 ( .A1(D[20]), .A2(n131), .ZN(n61) );
  OAI21_X1 U60 ( .B1(net55858), .B2(n135), .A(n62), .ZN(n11) );
  NAND2_X1 U61 ( .A1(D[21]), .A2(n131), .ZN(n62) );
  OAI21_X1 U62 ( .B1(net55859), .B2(n135), .A(n63), .ZN(n10) );
  NAND2_X1 U63 ( .A1(D[22]), .A2(n131), .ZN(n63) );
  OAI21_X1 U64 ( .B1(net55868), .B2(n135), .A(n64), .ZN(n1) );
  NAND2_X1 U65 ( .A1(D[31]), .A2(n131), .ZN(n64) );
  OAI21_X1 U66 ( .B1(net55842), .B2(n134), .A(n45), .ZN(n27) );
  NAND2_X1 U67 ( .A1(D[5]), .A2(n133), .ZN(n45) );
  OAI21_X1 U68 ( .B1(net55843), .B2(n134), .A(n46), .ZN(n26) );
  NAND2_X1 U69 ( .A1(D[6]), .A2(n133), .ZN(n46) );
  OAI21_X1 U70 ( .B1(net55845), .B2(n134), .A(n48), .ZN(n24) );
  NAND2_X1 U71 ( .A1(D[8]), .A2(n133), .ZN(n48) );
  OAI21_X1 U72 ( .B1(net55846), .B2(n134), .A(n49), .ZN(n23) );
  NAND2_X1 U73 ( .A1(D[9]), .A2(n133), .ZN(n49) );
  BUF_X1 U74 ( .A(ENABLE), .Z(n130) );
  BUF_X1 U75 ( .A(n85), .Z(n137) );
  BUF_X1 U76 ( .A(n85), .Z(n136) );
  BUF_X1 U77 ( .A(n85), .Z(n138) );
  MUX2_X1 U78 ( .A(Q[2]), .B(D[2]), .S(n135), .Z(n30) );
  MUX2_X1 U79 ( .A(n139), .B(D[0]), .S(n135), .Z(n32) );
  MUX2_X1 U80 ( .A(n119), .B(D[1]), .S(n135), .Z(n31) );
endmodule


module D_Reg_generic_N32_9 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55837, net55838, net55839, net55840, net55841, net55842,
         net55843, net55844, net55845, net55846, net55847, net55848, net55849,
         net55850, net55851, net55852, net55853, net55854, net55855, net55856,
         net55857, net55858, net55859, net55860, net55861, net55862, net55863,
         net55864, net55865, net55866, net55867, net55868, n73, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n106, n107, n108, n109, n110, n111, n112, n113, n114;
  assign n73 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n114), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n112), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n114), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n112), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n114), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n112), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n112), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n112), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n114), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n112), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n112), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n112), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n114), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n113), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n113), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n113), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n112), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n113), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n113), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n113), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n113), .Q(Q[11]), .QN(net55848)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n113), .Q(Q[10]), .QN(net55847)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n114), .Q(Q[9]), .QN(net55846)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n112), .Q(Q[8]), .QN(net55845)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n114), .Q(Q[7]), .QN(net55844)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n112), .Q(Q[6]), .QN(net55843)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n113), .Q(Q[5]), .QN(net55842)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n112), .Q(Q[4]), .QN(net55841)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n113), .Q(Q[3]), .QN(net55840)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n113), .Q(Q[2]), .QN(net55839)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n113), .Q(Q[1]), .QN(net55838)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n114), .Q(Q[0]), .QN(net55837)
         );
  BUF_X1 U2 ( .A(ENABLE), .Z(n107) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n106) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n108) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n110) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n109) );
  OAI21_X1 U7 ( .B1(net55838), .B2(n108), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(D[1]), .A2(n107), .ZN(n40) );
  OAI21_X1 U9 ( .B1(net55861), .B2(n108), .A(n34), .ZN(n8) );
  NAND2_X1 U10 ( .A1(D[24]), .A2(n106), .ZN(n34) );
  OAI21_X1 U11 ( .B1(net55862), .B2(n108), .A(n35), .ZN(n7) );
  NAND2_X1 U12 ( .A1(D[25]), .A2(n106), .ZN(n35) );
  OAI21_X1 U13 ( .B1(net55864), .B2(n108), .A(n37), .ZN(n5) );
  NAND2_X1 U14 ( .A1(D[27]), .A2(n106), .ZN(n37) );
  OAI21_X1 U15 ( .B1(net55865), .B2(n108), .A(n38), .ZN(n4) );
  NAND2_X1 U16 ( .A1(D[28]), .A2(n107), .ZN(n38) );
  OAI21_X1 U17 ( .B1(net55837), .B2(n109), .A(n39), .ZN(n32) );
  NAND2_X1 U18 ( .A1(D[0]), .A2(n107), .ZN(n39) );
  OAI21_X1 U19 ( .B1(net55839), .B2(n109), .A(n41), .ZN(n30) );
  NAND2_X1 U20 ( .A1(D[2]), .A2(n107), .ZN(n41) );
  OAI21_X1 U21 ( .B1(net55840), .B2(n109), .A(n43), .ZN(n29) );
  NAND2_X1 U22 ( .A1(D[3]), .A2(n107), .ZN(n43) );
  OAI21_X1 U23 ( .B1(net55847), .B2(n110), .A(n50), .ZN(n22) );
  NAND2_X1 U24 ( .A1(D[10]), .A2(n107), .ZN(n50) );
  OAI21_X1 U25 ( .B1(net55848), .B2(n110), .A(n51), .ZN(n21) );
  NAND2_X1 U26 ( .A1(D[11]), .A2(n107), .ZN(n51) );
  OAI21_X1 U27 ( .B1(net55849), .B2(n110), .A(n52), .ZN(n20) );
  NAND2_X1 U28 ( .A1(D[12]), .A2(n107), .ZN(n52) );
  OAI21_X1 U29 ( .B1(net55850), .B2(n110), .A(n54), .ZN(n19) );
  NAND2_X1 U30 ( .A1(D[13]), .A2(n107), .ZN(n54) );
  OAI21_X1 U31 ( .B1(net55851), .B2(n110), .A(n55), .ZN(n18) );
  NAND2_X1 U32 ( .A1(D[14]), .A2(n107), .ZN(n55) );
  OAI21_X1 U33 ( .B1(net55852), .B2(n110), .A(n56), .ZN(n17) );
  NAND2_X1 U34 ( .A1(D[15]), .A2(n107), .ZN(n56) );
  OAI21_X1 U35 ( .B1(net55853), .B2(n110), .A(n57), .ZN(n16) );
  NAND2_X1 U36 ( .A1(D[16]), .A2(n106), .ZN(n57) );
  OAI21_X1 U37 ( .B1(net55854), .B2(n110), .A(n58), .ZN(n15) );
  NAND2_X1 U38 ( .A1(D[17]), .A2(n106), .ZN(n58) );
  OAI21_X1 U39 ( .B1(net55855), .B2(n110), .A(n59), .ZN(n14) );
  NAND2_X1 U40 ( .A1(D[18]), .A2(n106), .ZN(n59) );
  OAI21_X1 U41 ( .B1(net55856), .B2(n110), .A(n60), .ZN(n13) );
  NAND2_X1 U42 ( .A1(D[19]), .A2(n106), .ZN(n60) );
  OAI21_X1 U43 ( .B1(net55863), .B2(n109), .A(n36), .ZN(n6) );
  NAND2_X1 U44 ( .A1(D[26]), .A2(n106), .ZN(n36) );
  OAI21_X1 U45 ( .B1(net55867), .B2(n110), .A(n53), .ZN(n2) );
  NAND2_X1 U46 ( .A1(D[30]), .A2(n107), .ZN(n53) );
  OAI21_X1 U47 ( .B1(net55868), .B2(n109), .A(n64), .ZN(n1) );
  NAND2_X1 U48 ( .A1(D[31]), .A2(n106), .ZN(n64) );
  OAI21_X1 U49 ( .B1(net55857), .B2(n111), .A(n61), .ZN(n12) );
  NAND2_X1 U50 ( .A1(D[20]), .A2(n106), .ZN(n61) );
  OAI21_X1 U51 ( .B1(net55858), .B2(n111), .A(n62), .ZN(n11) );
  NAND2_X1 U52 ( .A1(D[21]), .A2(n106), .ZN(n62) );
  OAI21_X1 U53 ( .B1(net55859), .B2(n111), .A(n63), .ZN(n10) );
  NAND2_X1 U54 ( .A1(D[22]), .A2(n106), .ZN(n63) );
  OAI21_X1 U55 ( .B1(net55841), .B2(n109), .A(n44), .ZN(n28) );
  NAND2_X1 U56 ( .A1(D[4]), .A2(n108), .ZN(n44) );
  OAI21_X1 U57 ( .B1(net55842), .B2(n109), .A(n45), .ZN(n27) );
  NAND2_X1 U58 ( .A1(D[5]), .A2(n108), .ZN(n45) );
  OAI21_X1 U59 ( .B1(net55843), .B2(n109), .A(n46), .ZN(n26) );
  NAND2_X1 U60 ( .A1(D[6]), .A2(n108), .ZN(n46) );
  OAI21_X1 U61 ( .B1(net55844), .B2(n109), .A(n47), .ZN(n25) );
  NAND2_X1 U62 ( .A1(D[7]), .A2(n108), .ZN(n47) );
  OAI21_X1 U63 ( .B1(net55845), .B2(n109), .A(n48), .ZN(n24) );
  NAND2_X1 U64 ( .A1(D[8]), .A2(n108), .ZN(n48) );
  OAI21_X1 U65 ( .B1(net55846), .B2(n110), .A(n49), .ZN(n23) );
  NAND2_X1 U66 ( .A1(D[9]), .A2(n108), .ZN(n49) );
  OAI21_X1 U67 ( .B1(net55866), .B2(n109), .A(n42), .ZN(n3) );
  NAND2_X1 U68 ( .A1(D[29]), .A2(n108), .ZN(n42) );
  OAI21_X1 U69 ( .B1(net55860), .B2(n109), .A(n33), .ZN(n9) );
  NAND2_X1 U70 ( .A1(n111), .A2(D[23]), .ZN(n33) );
  BUF_X1 U71 ( .A(n73), .Z(n113) );
  BUF_X1 U72 ( .A(n73), .Z(n112) );
  BUF_X1 U73 ( .A(n73), .Z(n114) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n111) );
endmodule


module mux41_generic_N32_0 ( A, B, C, D, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] S;
  output [31:0] Y;

  wire   [31:0] ABto2;
  wire   [31:0] CDto2;

  MUX21_GENERIC_N32_0 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_GENERIC_N32_19 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_GENERIC_N32_18 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(Y) );
endmodule


module mux41_generic_N5 ( A, B, C, D, S, Y );
  input [4:0] A;
  input [4:0] B;
  input [4:0] C;
  input [4:0] D;
  input [1:0] S;
  output [4:0] Y;

  wire   [4:0] ABto2;
  wire   [4:0] CDto2;

  MUX21_GENERIC_N5_0 M11 ( .A(A), .B(B), .S(S[0]), .Y(ABto2) );
  MUX21_GENERIC_N5_2 M12 ( .A(C), .B(D), .S(S[0]), .Y(CDto2) );
  MUX21_GENERIC_N5_1 M21 ( .A(ABto2), .B(CDto2), .S(S[1]), .Y(Y) );
endmodule


module register_file_gen_Nbit32_Nreg32 ( RESET, ENABLE, WR, RD1, RD2, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input RESET, ENABLE, WR, RD1, RD2;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N4403, N4405, N4407, N4409, N4411, N4413, N4415,
         N4417, N4419, N4421, N4423, N4425, N4427, N4429, N4431, N4433, N4435,
         N4437, N4439, N4441, N4443, N4445, N4447, N4449, N4451, N4453, N4455,
         N4457, N4459, N4461, N4463, N4465, N4467, N4469, N4471, N4473, N4475,
         N4477, N4479, N4481, N4483, N4485, N4487, N4489, N4491, N4493, N4495,
         N4497, N4499, N4501, N4503, N4505, N4507, N4509, N4511, N4513, N4515,
         N4517, N4519, N4521, N4523, N4525, N4527, N4529, n2500, n2503, n2506,
         n2509, n2512, n2515, n2518, n2521, n2524, n2527, n2530, n2533, n2536,
         n2539, n2542, n2545, n2548, n2551, n2554, n2557, n2560, n2563, n2566,
         n2569, n2572, n2575, n2578, n2581, n2584, n2587, n2590, n2593, n2596,
         n2599, n2602, n2605, n2608, n2611, n2614, n2617, n2620, n2623, n2626,
         n2629, n2632, n2635, n2638, n2641, n2644, n2647, n2650, n2653, n2656,
         n2659, n2662, n2665, n2668, n2671, n2674, n2677, n2680, n2683, n2686,
         n2689, n2692, n2695, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099;

  DLH_X1 \REGISTERS_reg[0][31]  ( .G(n3083), .D(n3084), .Q(\REGISTERS[0][31] )
         );
  DLH_X1 \REGISTERS_reg[0][30]  ( .G(n3081), .D(n3078), .Q(\REGISTERS[0][30] )
         );
  DLH_X1 \REGISTERS_reg[0][29]  ( .G(n3083), .D(n3075), .Q(\REGISTERS[0][29] )
         );
  DLH_X1 \REGISTERS_reg[0][28]  ( .G(n3081), .D(n3072), .Q(\REGISTERS[0][28] )
         );
  DLH_X1 \REGISTERS_reg[0][27]  ( .G(n3083), .D(n3069), .Q(\REGISTERS[0][27] )
         );
  DLH_X1 \REGISTERS_reg[0][26]  ( .G(n3081), .D(n3066), .Q(\REGISTERS[0][26] )
         );
  DLH_X1 \REGISTERS_reg[0][25]  ( .G(n3081), .D(n3063), .Q(\REGISTERS[0][25] )
         );
  DLH_X1 \REGISTERS_reg[0][24]  ( .G(n3081), .D(n3060), .Q(\REGISTERS[0][24] )
         );
  DLH_X1 \REGISTERS_reg[0][23]  ( .G(n3083), .D(n3057), .Q(\REGISTERS[0][23] )
         );
  DLH_X1 \REGISTERS_reg[0][22]  ( .G(n3081), .D(n3054), .Q(\REGISTERS[0][22] )
         );
  DLH_X1 \REGISTERS_reg[0][21]  ( .G(n3081), .D(n3051), .Q(\REGISTERS[0][21] )
         );
  DLH_X1 \REGISTERS_reg[0][20]  ( .G(n3082), .D(n3048), .Q(\REGISTERS[0][20] )
         );
  DLH_X1 \REGISTERS_reg[0][19]  ( .G(n3083), .D(n3045), .Q(\REGISTERS[0][19] )
         );
  DLH_X1 \REGISTERS_reg[0][18]  ( .G(n3082), .D(n3042), .Q(\REGISTERS[0][18] )
         );
  DLH_X1 \REGISTERS_reg[0][17]  ( .G(n3082), .D(n3039), .Q(\REGISTERS[0][17] )
         );
  DLH_X1 \REGISTERS_reg[0][16]  ( .G(n3082), .D(n3036), .Q(\REGISTERS[0][16] )
         );
  DLH_X1 \REGISTERS_reg[0][15]  ( .G(n3081), .D(n3033), .Q(\REGISTERS[0][15] )
         );
  DLH_X1 \REGISTERS_reg[0][14]  ( .G(n3082), .D(n3030), .Q(\REGISTERS[0][14] )
         );
  DLH_X1 \REGISTERS_reg[0][13]  ( .G(n3082), .D(n3027), .Q(\REGISTERS[0][13] )
         );
  DLH_X1 \REGISTERS_reg[0][12]  ( .G(n3082), .D(n3024), .Q(\REGISTERS[0][12] )
         );
  DLH_X1 \REGISTERS_reg[0][11]  ( .G(n3083), .D(n3021), .Q(\REGISTERS[0][11] )
         );
  DLH_X1 \REGISTERS_reg[0][10]  ( .G(n3083), .D(n3018), .Q(\REGISTERS[0][10] )
         );
  DLH_X1 \REGISTERS_reg[0][9]  ( .G(n3083), .D(n3015), .Q(\REGISTERS[0][9] )
         );
  DLH_X1 \REGISTERS_reg[0][8]  ( .G(n3081), .D(n3012), .Q(\REGISTERS[0][8] )
         );
  DLH_X1 \REGISTERS_reg[0][7]  ( .G(n3083), .D(n3009), .Q(\REGISTERS[0][7] )
         );
  DLH_X1 \REGISTERS_reg[0][6]  ( .G(n3081), .D(n3006), .Q(\REGISTERS[0][6] )
         );
  DLH_X1 \REGISTERS_reg[0][5]  ( .G(n3082), .D(n3003), .Q(\REGISTERS[0][5] )
         );
  DLH_X1 \REGISTERS_reg[0][4]  ( .G(n3081), .D(n3000), .Q(\REGISTERS[0][4] )
         );
  DLH_X1 \REGISTERS_reg[0][3]  ( .G(n3082), .D(n2997), .Q(\REGISTERS[0][3] )
         );
  DLH_X1 \REGISTERS_reg[0][2]  ( .G(n3082), .D(n2994), .Q(\REGISTERS[0][2] )
         );
  DLH_X1 \REGISTERS_reg[0][1]  ( .G(n3082), .D(n2991), .Q(\REGISTERS[0][1] )
         );
  DLH_X1 \REGISTERS_reg[0][0]  ( .G(n3083), .D(n2988), .Q(\REGISTERS[0][0] )
         );
  DLH_X1 \REGISTERS_reg[1][31]  ( .G(n2987), .D(n3085), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(n2985), .D(n3079), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(n2987), .D(n3076), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(n2985), .D(n3073), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(n2987), .D(n3070), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(n2985), .D(n3067), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(n2985), .D(n3064), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(n2985), .D(n3061), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(n2987), .D(n3058), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(n2985), .D(n3055), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(n2985), .D(n3052), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n2986), .D(n3049), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n2987), .D(n3046), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(n2986), .D(n3043), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(n2986), .D(n3040), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(n2986), .D(n3037), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(n2985), .D(n3034), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(n2986), .D(n3031), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(n2986), .D(n3028), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(n2986), .D(n3025), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n2987), .D(n3022), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(n2987), .D(n3019), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(n2987), .D(n3016), .Q(\REGISTERS[1][9] )
         );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(n2985), .D(n3013), .Q(\REGISTERS[1][8] )
         );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n2987), .D(n3010), .Q(\REGISTERS[1][7] )
         );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(n2985), .D(n3007), .Q(\REGISTERS[1][6] )
         );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n2986), .D(n3004), .Q(\REGISTERS[1][5] )
         );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(n2985), .D(n3001), .Q(\REGISTERS[1][4] )
         );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(n2986), .D(n2998), .Q(\REGISTERS[1][3] )
         );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(n2986), .D(n2995), .Q(\REGISTERS[1][2] )
         );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(n2986), .D(n2992), .Q(\REGISTERS[1][1] )
         );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n2987), .D(n2989), .Q(\REGISTERS[1][0] )
         );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(n2984), .D(n3085), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(n2982), .D(n3079), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(n2984), .D(n3076), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(n2982), .D(n3073), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(n2984), .D(n3070), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(n2982), .D(n3067), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(n2982), .D(n3064), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(n2982), .D(n3061), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n2984), .D(n3058), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n2982), .D(n3055), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(n2982), .D(n3052), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(n2983), .D(n3049), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n2984), .D(n3046), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(n2983), .D(n3043), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n2983), .D(n3040), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(n2983), .D(n3037), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(n2982), .D(n3034), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(n2983), .D(n3031), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(n2983), .D(n3028), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(n2983), .D(n3025), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(n2984), .D(n3022), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n2984), .D(n3019), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(n2984), .D(n3016), .Q(\REGISTERS[2][9] )
         );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(n2982), .D(n3013), .Q(\REGISTERS[2][8] )
         );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n2984), .D(n3010), .Q(\REGISTERS[2][7] )
         );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(n2982), .D(n3007), .Q(\REGISTERS[2][6] )
         );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(n2983), .D(n3004), .Q(\REGISTERS[2][5] )
         );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(n2982), .D(n3001), .Q(\REGISTERS[2][4] )
         );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(n2983), .D(n2998), .Q(\REGISTERS[2][3] )
         );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(n2983), .D(n2995), .Q(\REGISTERS[2][2] )
         );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(n2983), .D(n2992), .Q(\REGISTERS[2][1] )
         );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(n2984), .D(n2989), .Q(\REGISTERS[2][0] )
         );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(n2981), .D(n3085), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(n2979), .D(n3079), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(n2981), .D(n3076), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(n2979), .D(n3073), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(n2981), .D(n3070), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(n2979), .D(n3067), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(n2979), .D(n3064), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(n2979), .D(n3061), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n2981), .D(n3058), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n2979), .D(n3055), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(n2979), .D(n3052), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(n2980), .D(n3049), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n2981), .D(n3046), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(n2980), .D(n3043), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n2980), .D(n3040), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(n2980), .D(n3037), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(n2979), .D(n3034), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(n2980), .D(n3031), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(n2980), .D(n3028), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(n2980), .D(n3025), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(n2981), .D(n3022), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n2981), .D(n3019), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(n2981), .D(n3016), .Q(\REGISTERS[3][9] )
         );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(n2979), .D(n3013), .Q(\REGISTERS[3][8] )
         );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n2981), .D(n3010), .Q(\REGISTERS[3][7] )
         );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(n2979), .D(n3007), .Q(\REGISTERS[3][6] )
         );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(n2980), .D(n3004), .Q(\REGISTERS[3][5] )
         );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(n2979), .D(n3001), .Q(\REGISTERS[3][4] )
         );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(n2980), .D(n2998), .Q(\REGISTERS[3][3] )
         );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(n2980), .D(n2995), .Q(\REGISTERS[3][2] )
         );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(n2980), .D(n2992), .Q(\REGISTERS[3][1] )
         );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(n2981), .D(n2989), .Q(\REGISTERS[3][0] )
         );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(n2978), .D(n3085), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(n2976), .D(n3079), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(n2978), .D(n3076), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(n2976), .D(n3073), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(n2978), .D(n3070), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(n2976), .D(n3067), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(n2976), .D(n3064), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(n2976), .D(n3061), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n2978), .D(n3058), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n2976), .D(n3055), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(n2976), .D(n3052), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(n2977), .D(n3049), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n2978), .D(n3046), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(n2977), .D(n3043), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n2977), .D(n3040), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(n2977), .D(n3037), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(n2976), .D(n3034), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(n2977), .D(n3031), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(n2977), .D(n3028), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(n2977), .D(n3025), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(n2978), .D(n3022), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n2978), .D(n3019), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(n2978), .D(n3016), .Q(\REGISTERS[4][9] )
         );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(n2976), .D(n3013), .Q(\REGISTERS[4][8] )
         );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(n2978), .D(n3010), .Q(\REGISTERS[4][7] )
         );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(n2976), .D(n3007), .Q(\REGISTERS[4][6] )
         );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(n2977), .D(n3004), .Q(\REGISTERS[4][5] )
         );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(n2976), .D(n3001), .Q(\REGISTERS[4][4] )
         );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(n2977), .D(n2998), .Q(\REGISTERS[4][3] )
         );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(n2977), .D(n2995), .Q(\REGISTERS[4][2] )
         );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(n2977), .D(n2992), .Q(\REGISTERS[4][1] )
         );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n2978), .D(n2989), .Q(\REGISTERS[4][0] )
         );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(n2975), .D(n3085), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(n2973), .D(n3079), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(n2975), .D(n3076), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(n2973), .D(n3073), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(n2975), .D(n3070), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(n2973), .D(n3067), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(n2973), .D(n3064), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(n2973), .D(n3061), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n2975), .D(n3058), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n2973), .D(n3055), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(n2973), .D(n3052), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(n2974), .D(n3049), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n2975), .D(n3046), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(n2974), .D(n3043), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n2974), .D(n3040), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(n2974), .D(n3037), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(n2973), .D(n3034), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(n2974), .D(n3031), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(n2974), .D(n3028), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(n2974), .D(n3025), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(n2975), .D(n3022), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n2975), .D(n3019), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(n2975), .D(n3016), .Q(\REGISTERS[5][9] )
         );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(n2973), .D(n3013), .Q(\REGISTERS[5][8] )
         );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n2975), .D(n3010), .Q(\REGISTERS[5][7] )
         );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(n2973), .D(n3007), .Q(\REGISTERS[5][6] )
         );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(n2974), .D(n3004), .Q(\REGISTERS[5][5] )
         );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(n2973), .D(n3001), .Q(\REGISTERS[5][4] )
         );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(n2974), .D(n2998), .Q(\REGISTERS[5][3] )
         );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(n2974), .D(n2995), .Q(\REGISTERS[5][2] )
         );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(n2974), .D(n2992), .Q(\REGISTERS[5][1] )
         );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(n2975), .D(n2989), .Q(\REGISTERS[5][0] )
         );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(n2972), .D(n3085), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(n2970), .D(n3079), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(n2972), .D(n3076), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(n2970), .D(n3073), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(n2972), .D(n3070), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(n2970), .D(n3067), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(n2970), .D(n3064), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(n2970), .D(n3061), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n2972), .D(n3058), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n2970), .D(n3055), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(n2970), .D(n3052), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(n2971), .D(n3049), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n2972), .D(n3046), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(n2971), .D(n3043), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n2971), .D(n3040), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(n2971), .D(n3037), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(n2970), .D(n3034), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(n2971), .D(n3031), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(n2971), .D(n3028), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(n2971), .D(n3025), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(n2972), .D(n3022), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n2972), .D(n3019), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(n2972), .D(n3016), .Q(\REGISTERS[6][9] )
         );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(n2970), .D(n3013), .Q(\REGISTERS[6][8] )
         );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(n2972), .D(n3010), .Q(\REGISTERS[6][7] )
         );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(n2970), .D(n3007), .Q(\REGISTERS[6][6] )
         );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(n2971), .D(n3004), .Q(\REGISTERS[6][5] )
         );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(n2970), .D(n3001), .Q(\REGISTERS[6][4] )
         );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(n2971), .D(n2998), .Q(\REGISTERS[6][3] )
         );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(n2971), .D(n2995), .Q(\REGISTERS[6][2] )
         );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(n2971), .D(n2992), .Q(\REGISTERS[6][1] )
         );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n2972), .D(n2989), .Q(\REGISTERS[6][0] )
         );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(n2969), .D(n3085), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(n2967), .D(n3079), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(n2969), .D(n3076), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(n2967), .D(n3073), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(n2969), .D(n3070), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(n2967), .D(n3067), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(n2967), .D(n3064), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(n2967), .D(n3061), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n2969), .D(n3058), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n2967), .D(n3055), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(n2967), .D(n3052), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(n2968), .D(n3049), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n2969), .D(n3046), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(n2968), .D(n3043), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n2968), .D(n3040), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(n2968), .D(n3037), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(n2967), .D(n3034), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(n2968), .D(n3031), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(n2968), .D(n3028), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(n2968), .D(n3025), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(n2969), .D(n3022), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n2969), .D(n3019), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(n2969), .D(n3016), .Q(\REGISTERS[7][9] )
         );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(n2967), .D(n3013), .Q(\REGISTERS[7][8] )
         );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n2969), .D(n3010), .Q(\REGISTERS[7][7] )
         );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(n2967), .D(n3007), .Q(\REGISTERS[7][6] )
         );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(n2968), .D(n3004), .Q(\REGISTERS[7][5] )
         );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(n2967), .D(n3001), .Q(\REGISTERS[7][4] )
         );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(n2968), .D(n2998), .Q(\REGISTERS[7][3] )
         );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(n2968), .D(n2995), .Q(\REGISTERS[7][2] )
         );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(n2968), .D(n2992), .Q(\REGISTERS[7][1] )
         );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(n2969), .D(n2989), .Q(\REGISTERS[7][0] )
         );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(n2966), .D(n3085), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(n2964), .D(n3079), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(n2966), .D(n3076), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(n2964), .D(n3073), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(n2966), .D(n3070), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(n2964), .D(n3067), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(n2964), .D(n3064), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(n2964), .D(n3061), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n2966), .D(n3058), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n2964), .D(n3055), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(n2964), .D(n3052), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(n2965), .D(n3049), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n2966), .D(n3046), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(n2965), .D(n3043), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n2965), .D(n3040), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(n2965), .D(n3037), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(n2964), .D(n3034), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(n2965), .D(n3031), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(n2965), .D(n3028), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(n2965), .D(n3025), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(n2966), .D(n3022), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n2966), .D(n3019), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(n2966), .D(n3016), .Q(\REGISTERS[8][9] )
         );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(n2964), .D(n3013), .Q(\REGISTERS[8][8] )
         );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n2966), .D(n3010), .Q(\REGISTERS[8][7] )
         );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(n2964), .D(n3007), .Q(\REGISTERS[8][6] )
         );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(n2965), .D(n3004), .Q(\REGISTERS[8][5] )
         );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(n2964), .D(n3001), .Q(\REGISTERS[8][4] )
         );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(n2965), .D(n2998), .Q(\REGISTERS[8][3] )
         );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(n2965), .D(n2995), .Q(\REGISTERS[8][2] )
         );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(n2965), .D(n2992), .Q(\REGISTERS[8][1] )
         );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(n2966), .D(n2989), .Q(\REGISTERS[8][0] )
         );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(n2963), .D(n3085), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(n2961), .D(n3079), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(n2963), .D(n3076), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(n2961), .D(n3073), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(n2963), .D(n3070), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(n2961), .D(n3067), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(n2961), .D(n3064), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(n2961), .D(n3061), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n2963), .D(n3058), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n2961), .D(n3055), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(n2961), .D(n3052), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(n2962), .D(n3049), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n2963), .D(n3046), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(n2962), .D(n3043), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n2962), .D(n3040), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(n2962), .D(n3037), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(n2961), .D(n3034), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(n2962), .D(n3031), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(n2962), .D(n3028), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(n2962), .D(n3025), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(n2963), .D(n3022), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n2963), .D(n3019), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(n2963), .D(n3016), .Q(\REGISTERS[9][9] )
         );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(n2961), .D(n3013), .Q(\REGISTERS[9][8] )
         );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n2963), .D(n3010), .Q(\REGISTERS[9][7] )
         );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(n2961), .D(n3007), .Q(\REGISTERS[9][6] )
         );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(n2962), .D(n3004), .Q(\REGISTERS[9][5] )
         );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(n2961), .D(n3001), .Q(\REGISTERS[9][4] )
         );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(n2962), .D(n2998), .Q(\REGISTERS[9][3] )
         );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(n2962), .D(n2995), .Q(\REGISTERS[9][2] )
         );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(n2962), .D(n2992), .Q(\REGISTERS[9][1] )
         );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(n2963), .D(n2989), .Q(\REGISTERS[9][0] )
         );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(n2960), .D(n3085), .Q(
        \REGISTERS[10][31] ) );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(n2958), .D(n3079), .Q(
        \REGISTERS[10][30] ) );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(n2960), .D(n3076), .Q(
        \REGISTERS[10][29] ) );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(n2958), .D(n3073), .Q(
        \REGISTERS[10][28] ) );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(n2960), .D(n3070), .Q(
        \REGISTERS[10][27] ) );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(n2958), .D(n3067), .Q(
        \REGISTERS[10][26] ) );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(n2958), .D(n3064), .Q(
        \REGISTERS[10][25] ) );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(n2958), .D(n3061), .Q(
        \REGISTERS[10][24] ) );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n2960), .D(n3058), .Q(
        \REGISTERS[10][23] ) );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(n2958), .D(n3055), .Q(
        \REGISTERS[10][22] ) );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(n2958), .D(n3052), .Q(
        \REGISTERS[10][21] ) );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(n2959), .D(n3049), .Q(
        \REGISTERS[10][20] ) );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n2960), .D(n3046), .Q(
        \REGISTERS[10][19] ) );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(n2959), .D(n3043), .Q(
        \REGISTERS[10][18] ) );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(n2959), .D(n3040), .Q(
        \REGISTERS[10][17] ) );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n2959), .D(n3037), .Q(
        \REGISTERS[10][16] ) );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(n2958), .D(n3034), .Q(
        \REGISTERS[10][15] ) );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(n2959), .D(n3031), .Q(
        \REGISTERS[10][14] ) );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n2959), .D(n3028), .Q(
        \REGISTERS[10][13] ) );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(n2959), .D(n3025), .Q(
        \REGISTERS[10][12] ) );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n2960), .D(n3022), .Q(
        \REGISTERS[10][11] ) );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n2960), .D(n3019), .Q(
        \REGISTERS[10][10] ) );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(n2960), .D(n3016), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(n2958), .D(n3013), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(n2960), .D(n3010), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(n2958), .D(n3007), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(n2959), .D(n3004), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(n2958), .D(n3001), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(n2959), .D(n2998), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(n2959), .D(n2995), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(n2959), .D(n2992), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(n2960), .D(n2989), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(n2957), .D(n3086), .Q(
        \REGISTERS[11][31] ) );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(n2955), .D(n3080), .Q(
        \REGISTERS[11][30] ) );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(n2957), .D(n3077), .Q(
        \REGISTERS[11][29] ) );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(n2955), .D(n3074), .Q(
        \REGISTERS[11][28] ) );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(n2957), .D(n3071), .Q(
        \REGISTERS[11][27] ) );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(n2955), .D(n3068), .Q(
        \REGISTERS[11][26] ) );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(n2955), .D(n3065), .Q(
        \REGISTERS[11][25] ) );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(n2955), .D(n3062), .Q(
        \REGISTERS[11][24] ) );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n2957), .D(n3059), .Q(
        \REGISTERS[11][23] ) );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n2955), .D(n3056), .Q(
        \REGISTERS[11][22] ) );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(n2955), .D(n3053), .Q(
        \REGISTERS[11][21] ) );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(n2956), .D(n3050), .Q(
        \REGISTERS[11][20] ) );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n2957), .D(n3047), .Q(
        \REGISTERS[11][19] ) );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(n2956), .D(n3044), .Q(
        \REGISTERS[11][18] ) );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n2956), .D(n3041), .Q(
        \REGISTERS[11][17] ) );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(n2956), .D(n3038), .Q(
        \REGISTERS[11][16] ) );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(n2955), .D(n3035), .Q(
        \REGISTERS[11][15] ) );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(n2956), .D(n3032), .Q(
        \REGISTERS[11][14] ) );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(n2956), .D(n3029), .Q(
        \REGISTERS[11][13] ) );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(n2956), .D(n3026), .Q(
        \REGISTERS[11][12] ) );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(n2957), .D(n3023), .Q(
        \REGISTERS[11][11] ) );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n2957), .D(n3020), .Q(
        \REGISTERS[11][10] ) );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(n2957), .D(n3017), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(n2955), .D(n3014), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n2957), .D(n3011), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(n2955), .D(n3008), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(n2956), .D(n3005), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(n2955), .D(n3002), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(n2956), .D(n2999), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(n2956), .D(n2996), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(n2956), .D(n2993), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(n2957), .D(n2990), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(n2954), .D(n3086), .Q(
        \REGISTERS[12][31] ) );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(n2952), .D(n3080), .Q(
        \REGISTERS[12][30] ) );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(n2954), .D(n3077), .Q(
        \REGISTERS[12][29] ) );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(n2952), .D(n3074), .Q(
        \REGISTERS[12][28] ) );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(n2954), .D(n3071), .Q(
        \REGISTERS[12][27] ) );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(n2952), .D(n3068), .Q(
        \REGISTERS[12][26] ) );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(n2952), .D(n3065), .Q(
        \REGISTERS[12][25] ) );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(n2952), .D(n3062), .Q(
        \REGISTERS[12][24] ) );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n2954), .D(n3059), .Q(
        \REGISTERS[12][23] ) );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n2952), .D(n3056), .Q(
        \REGISTERS[12][22] ) );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(n2952), .D(n3053), .Q(
        \REGISTERS[12][21] ) );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(n2953), .D(n3050), .Q(
        \REGISTERS[12][20] ) );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n2954), .D(n3047), .Q(
        \REGISTERS[12][19] ) );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(n2953), .D(n3044), .Q(
        \REGISTERS[12][18] ) );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n2953), .D(n3041), .Q(
        \REGISTERS[12][17] ) );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(n2953), .D(n3038), .Q(
        \REGISTERS[12][16] ) );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(n2952), .D(n3035), .Q(
        \REGISTERS[12][15] ) );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(n2953), .D(n3032), .Q(
        \REGISTERS[12][14] ) );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(n2953), .D(n3029), .Q(
        \REGISTERS[12][13] ) );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(n2953), .D(n3026), .Q(
        \REGISTERS[12][12] ) );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n2954), .D(n3023), .Q(
        \REGISTERS[12][11] ) );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n2954), .D(n3020), .Q(
        \REGISTERS[12][10] ) );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(n2954), .D(n3017), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(n2952), .D(n3014), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(n2954), .D(n3011), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(n2952), .D(n3008), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(n2953), .D(n3005), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(n2952), .D(n3002), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(n2953), .D(n2999), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(n2953), .D(n2996), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(n2953), .D(n2993), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(n2954), .D(n2990), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(n2951), .D(n3086), .Q(
        \REGISTERS[13][31] ) );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(n2949), .D(n3080), .Q(
        \REGISTERS[13][30] ) );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(n2951), .D(n3077), .Q(
        \REGISTERS[13][29] ) );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(n2949), .D(n3074), .Q(
        \REGISTERS[13][28] ) );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(n2951), .D(n3071), .Q(
        \REGISTERS[13][27] ) );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(n2949), .D(n3068), .Q(
        \REGISTERS[13][26] ) );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(n2949), .D(n3065), .Q(
        \REGISTERS[13][25] ) );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(n2949), .D(n3062), .Q(
        \REGISTERS[13][24] ) );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n2951), .D(n3059), .Q(
        \REGISTERS[13][23] ) );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n2949), .D(n3056), .Q(
        \REGISTERS[13][22] ) );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(n2949), .D(n3053), .Q(
        \REGISTERS[13][21] ) );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(n2950), .D(n3050), .Q(
        \REGISTERS[13][20] ) );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n2951), .D(n3047), .Q(
        \REGISTERS[13][19] ) );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(n2950), .D(n3044), .Q(
        \REGISTERS[13][18] ) );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n2950), .D(n3041), .Q(
        \REGISTERS[13][17] ) );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(n2950), .D(n3038), .Q(
        \REGISTERS[13][16] ) );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(n2949), .D(n3035), .Q(
        \REGISTERS[13][15] ) );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(n2950), .D(n3032), .Q(
        \REGISTERS[13][14] ) );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(n2950), .D(n3029), .Q(
        \REGISTERS[13][13] ) );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(n2950), .D(n3026), .Q(
        \REGISTERS[13][12] ) );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(n2951), .D(n3023), .Q(
        \REGISTERS[13][11] ) );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n2951), .D(n3020), .Q(
        \REGISTERS[13][10] ) );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(n2951), .D(n3017), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(n2949), .D(n3014), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n2951), .D(n3011), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(n2949), .D(n3008), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(n2950), .D(n3005), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(n2949), .D(n3002), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(n2950), .D(n2999), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(n2950), .D(n2996), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(n2950), .D(n2993), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(n2951), .D(n2990), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(n2948), .D(n3086), .Q(
        \REGISTERS[14][31] ) );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(n2946), .D(n3080), .Q(
        \REGISTERS[14][30] ) );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(n2948), .D(n3077), .Q(
        \REGISTERS[14][29] ) );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(n2946), .D(n3074), .Q(
        \REGISTERS[14][28] ) );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(n2948), .D(n3071), .Q(
        \REGISTERS[14][27] ) );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(n2946), .D(n3068), .Q(
        \REGISTERS[14][26] ) );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(n2946), .D(n3065), .Q(
        \REGISTERS[14][25] ) );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(n2946), .D(n3062), .Q(
        \REGISTERS[14][24] ) );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n2948), .D(n3059), .Q(
        \REGISTERS[14][23] ) );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n2946), .D(n3056), .Q(
        \REGISTERS[14][22] ) );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(n2946), .D(n3053), .Q(
        \REGISTERS[14][21] ) );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(n2947), .D(n3050), .Q(
        \REGISTERS[14][20] ) );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n2948), .D(n3047), .Q(
        \REGISTERS[14][19] ) );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(n2947), .D(n3044), .Q(
        \REGISTERS[14][18] ) );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n2947), .D(n3041), .Q(
        \REGISTERS[14][17] ) );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(n2947), .D(n3038), .Q(
        \REGISTERS[14][16] ) );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(n2946), .D(n3035), .Q(
        \REGISTERS[14][15] ) );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(n2947), .D(n3032), .Q(
        \REGISTERS[14][14] ) );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(n2947), .D(n3029), .Q(
        \REGISTERS[14][13] ) );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(n2947), .D(n3026), .Q(
        \REGISTERS[14][12] ) );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(n2948), .D(n3023), .Q(
        \REGISTERS[14][11] ) );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n2948), .D(n3020), .Q(
        \REGISTERS[14][10] ) );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(n2948), .D(n3017), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(n2946), .D(n3014), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n2948), .D(n3011), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(n2946), .D(n3008), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(n2947), .D(n3005), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(n2946), .D(n3002), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(n2947), .D(n2999), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(n2947), .D(n2996), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(n2947), .D(n2993), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(n2948), .D(n2990), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(n2945), .D(n3086), .Q(
        \REGISTERS[15][31] ) );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(n2943), .D(n3080), .Q(
        \REGISTERS[15][30] ) );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(n2945), .D(n3077), .Q(
        \REGISTERS[15][29] ) );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(n2943), .D(n3074), .Q(
        \REGISTERS[15][28] ) );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(n2945), .D(n3071), .Q(
        \REGISTERS[15][27] ) );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(n2943), .D(n3068), .Q(
        \REGISTERS[15][26] ) );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(n2943), .D(n3065), .Q(
        \REGISTERS[15][25] ) );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(n2943), .D(n3062), .Q(
        \REGISTERS[15][24] ) );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n2945), .D(n3059), .Q(
        \REGISTERS[15][23] ) );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n2943), .D(n3056), .Q(
        \REGISTERS[15][22] ) );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(n2943), .D(n3053), .Q(
        \REGISTERS[15][21] ) );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(n2944), .D(n3050), .Q(
        \REGISTERS[15][20] ) );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n2945), .D(n3047), .Q(
        \REGISTERS[15][19] ) );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(n2944), .D(n3044), .Q(
        \REGISTERS[15][18] ) );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n2944), .D(n3041), .Q(
        \REGISTERS[15][17] ) );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(n2944), .D(n3038), .Q(
        \REGISTERS[15][16] ) );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(n2943), .D(n3035), .Q(
        \REGISTERS[15][15] ) );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(n2944), .D(n3032), .Q(
        \REGISTERS[15][14] ) );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(n2944), .D(n3029), .Q(
        \REGISTERS[15][13] ) );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(n2944), .D(n3026), .Q(
        \REGISTERS[15][12] ) );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(n2945), .D(n3023), .Q(
        \REGISTERS[15][11] ) );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n2945), .D(n3020), .Q(
        \REGISTERS[15][10] ) );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(n2945), .D(n3017), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(n2943), .D(n3014), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n2945), .D(n3011), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(n2943), .D(n3008), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(n2944), .D(n3005), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(n2943), .D(n3002), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(n2944), .D(n2999), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(n2944), .D(n2996), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(n2944), .D(n2993), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(n2945), .D(n2990), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(n2942), .D(n3086), .Q(
        \REGISTERS[16][31] ) );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(n2940), .D(n3080), .Q(
        \REGISTERS[16][30] ) );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(n2942), .D(n3077), .Q(
        \REGISTERS[16][29] ) );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(n2940), .D(n3074), .Q(
        \REGISTERS[16][28] ) );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(n2942), .D(n3071), .Q(
        \REGISTERS[16][27] ) );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(n2940), .D(n3068), .Q(
        \REGISTERS[16][26] ) );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(n2940), .D(n3065), .Q(
        \REGISTERS[16][25] ) );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(n2940), .D(n3062), .Q(
        \REGISTERS[16][24] ) );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n2942), .D(n3059), .Q(
        \REGISTERS[16][23] ) );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n2940), .D(n3056), .Q(
        \REGISTERS[16][22] ) );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(n2940), .D(n3053), .Q(
        \REGISTERS[16][21] ) );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(n2941), .D(n3050), .Q(
        \REGISTERS[16][20] ) );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n2942), .D(n3047), .Q(
        \REGISTERS[16][19] ) );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(n2941), .D(n3044), .Q(
        \REGISTERS[16][18] ) );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n2941), .D(n3041), .Q(
        \REGISTERS[16][17] ) );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(n2941), .D(n3038), .Q(
        \REGISTERS[16][16] ) );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(n2940), .D(n3035), .Q(
        \REGISTERS[16][15] ) );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(n2941), .D(n3032), .Q(
        \REGISTERS[16][14] ) );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(n2941), .D(n3029), .Q(
        \REGISTERS[16][13] ) );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(n2941), .D(n3026), .Q(
        \REGISTERS[16][12] ) );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(n2942), .D(n3023), .Q(
        \REGISTERS[16][11] ) );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n2942), .D(n3020), .Q(
        \REGISTERS[16][10] ) );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(n2942), .D(n3017), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(n2940), .D(n3014), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n2942), .D(n3011), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(n2940), .D(n3008), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(n2941), .D(n3005), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(n2940), .D(n3002), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(n2941), .D(n2999), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(n2941), .D(n2996), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(n2941), .D(n2993), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(n2942), .D(n2990), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(n2939), .D(n3086), .Q(
        \REGISTERS[17][31] ) );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(n2937), .D(n3080), .Q(
        \REGISTERS[17][30] ) );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(n2939), .D(n3077), .Q(
        \REGISTERS[17][29] ) );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(n2937), .D(n3074), .Q(
        \REGISTERS[17][28] ) );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(n2939), .D(n3071), .Q(
        \REGISTERS[17][27] ) );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(n2937), .D(n3068), .Q(
        \REGISTERS[17][26] ) );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(n2937), .D(n3065), .Q(
        \REGISTERS[17][25] ) );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(n2937), .D(n3062), .Q(
        \REGISTERS[17][24] ) );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n2939), .D(n3059), .Q(
        \REGISTERS[17][23] ) );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n2937), .D(n3056), .Q(
        \REGISTERS[17][22] ) );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(n2937), .D(n3053), .Q(
        \REGISTERS[17][21] ) );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(n2938), .D(n3050), .Q(
        \REGISTERS[17][20] ) );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n2939), .D(n3047), .Q(
        \REGISTERS[17][19] ) );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(n2938), .D(n3044), .Q(
        \REGISTERS[17][18] ) );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n2938), .D(n3041), .Q(
        \REGISTERS[17][17] ) );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(n2938), .D(n3038), .Q(
        \REGISTERS[17][16] ) );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(n2937), .D(n3035), .Q(
        \REGISTERS[17][15] ) );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(n2938), .D(n3032), .Q(
        \REGISTERS[17][14] ) );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(n2938), .D(n3029), .Q(
        \REGISTERS[17][13] ) );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(n2938), .D(n3026), .Q(
        \REGISTERS[17][12] ) );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(n2939), .D(n3023), .Q(
        \REGISTERS[17][11] ) );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n2939), .D(n3020), .Q(
        \REGISTERS[17][10] ) );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(n2939), .D(n3017), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(n2937), .D(n3014), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n2939), .D(n3011), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(n2937), .D(n3008), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(n2938), .D(n3005), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(n2937), .D(n3002), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(n2938), .D(n2999), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(n2938), .D(n2996), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(n2938), .D(n2993), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(n2939), .D(n2990), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(n2936), .D(n3086), .Q(
        \REGISTERS[18][31] ) );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(n2934), .D(n3080), .Q(
        \REGISTERS[18][30] ) );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(n2936), .D(n3077), .Q(
        \REGISTERS[18][29] ) );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(n2934), .D(n3074), .Q(
        \REGISTERS[18][28] ) );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(n2936), .D(n3071), .Q(
        \REGISTERS[18][27] ) );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(n2934), .D(n3068), .Q(
        \REGISTERS[18][26] ) );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(n2934), .D(n3065), .Q(
        \REGISTERS[18][25] ) );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(n2934), .D(n3062), .Q(
        \REGISTERS[18][24] ) );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n2936), .D(n3059), .Q(
        \REGISTERS[18][23] ) );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n2934), .D(n3056), .Q(
        \REGISTERS[18][22] ) );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(n2934), .D(n3053), .Q(
        \REGISTERS[18][21] ) );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(n2935), .D(n3050), .Q(
        \REGISTERS[18][20] ) );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n2936), .D(n3047), .Q(
        \REGISTERS[18][19] ) );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(n2935), .D(n3044), .Q(
        \REGISTERS[18][18] ) );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n2935), .D(n3041), .Q(
        \REGISTERS[18][17] ) );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(n2935), .D(n3038), .Q(
        \REGISTERS[18][16] ) );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(n2934), .D(n3035), .Q(
        \REGISTERS[18][15] ) );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(n2935), .D(n3032), .Q(
        \REGISTERS[18][14] ) );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(n2935), .D(n3029), .Q(
        \REGISTERS[18][13] ) );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(n2935), .D(n3026), .Q(
        \REGISTERS[18][12] ) );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(n2936), .D(n3023), .Q(
        \REGISTERS[18][11] ) );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n2936), .D(n3020), .Q(
        \REGISTERS[18][10] ) );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(n2936), .D(n3017), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(n2934), .D(n3014), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n2936), .D(n3011), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(n2934), .D(n3008), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(n2935), .D(n3005), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(n2934), .D(n3002), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(n2935), .D(n2999), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(n2935), .D(n2996), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(n2935), .D(n2993), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(n2936), .D(n2990), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(n2933), .D(n3086), .Q(
        \REGISTERS[19][31] ) );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(n2931), .D(n3080), .Q(
        \REGISTERS[19][30] ) );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(n2933), .D(n3077), .Q(
        \REGISTERS[19][29] ) );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(n2931), .D(n3074), .Q(
        \REGISTERS[19][28] ) );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(n2933), .D(n3071), .Q(
        \REGISTERS[19][27] ) );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(n2931), .D(n3068), .Q(
        \REGISTERS[19][26] ) );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(n2931), .D(n3065), .Q(
        \REGISTERS[19][25] ) );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(n2931), .D(n3062), .Q(
        \REGISTERS[19][24] ) );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n2933), .D(n3059), .Q(
        \REGISTERS[19][23] ) );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n2931), .D(n3056), .Q(
        \REGISTERS[19][22] ) );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(n2931), .D(n3053), .Q(
        \REGISTERS[19][21] ) );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(n2932), .D(n3050), .Q(
        \REGISTERS[19][20] ) );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n2933), .D(n3047), .Q(
        \REGISTERS[19][19] ) );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(n2932), .D(n3044), .Q(
        \REGISTERS[19][18] ) );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n2932), .D(n3041), .Q(
        \REGISTERS[19][17] ) );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(n2932), .D(n3038), .Q(
        \REGISTERS[19][16] ) );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(n2931), .D(n3035), .Q(
        \REGISTERS[19][15] ) );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(n2932), .D(n3032), .Q(
        \REGISTERS[19][14] ) );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(n2932), .D(n3029), .Q(
        \REGISTERS[19][13] ) );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(n2932), .D(n3026), .Q(
        \REGISTERS[19][12] ) );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(n2933), .D(n3023), .Q(
        \REGISTERS[19][11] ) );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n2933), .D(n3020), .Q(
        \REGISTERS[19][10] ) );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(n2933), .D(n3017), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(n2931), .D(n3014), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n2933), .D(n3011), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(n2931), .D(n3008), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(n2932), .D(n3005), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(n2931), .D(n3002), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(n2932), .D(n2999), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(n2932), .D(n2996), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(n2932), .D(n2993), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(n2933), .D(n2990), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(n2930), .D(n3086), .Q(
        \REGISTERS[20][31] ) );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(n2928), .D(n3080), .Q(
        \REGISTERS[20][30] ) );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(n2930), .D(n3077), .Q(
        \REGISTERS[20][29] ) );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(n2928), .D(n3074), .Q(
        \REGISTERS[20][28] ) );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(n2930), .D(n3071), .Q(
        \REGISTERS[20][27] ) );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(n2928), .D(n3068), .Q(
        \REGISTERS[20][26] ) );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(n2928), .D(n3065), .Q(
        \REGISTERS[20][25] ) );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(n2928), .D(n3062), .Q(
        \REGISTERS[20][24] ) );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n2930), .D(n3059), .Q(
        \REGISTERS[20][23] ) );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n2928), .D(n3056), .Q(
        \REGISTERS[20][22] ) );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(n2928), .D(n3053), .Q(
        \REGISTERS[20][21] ) );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(n2929), .D(n3050), .Q(
        \REGISTERS[20][20] ) );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n2930), .D(n3047), .Q(
        \REGISTERS[20][19] ) );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(n2929), .D(n3044), .Q(
        \REGISTERS[20][18] ) );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n2929), .D(n3041), .Q(
        \REGISTERS[20][17] ) );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(n2929), .D(n3038), .Q(
        \REGISTERS[20][16] ) );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(n2928), .D(n3035), .Q(
        \REGISTERS[20][15] ) );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(n2929), .D(n3032), .Q(
        \REGISTERS[20][14] ) );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(n2929), .D(n3029), .Q(
        \REGISTERS[20][13] ) );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(n2929), .D(n3026), .Q(
        \REGISTERS[20][12] ) );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(n2930), .D(n3023), .Q(
        \REGISTERS[20][11] ) );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n2930), .D(n3020), .Q(
        \REGISTERS[20][10] ) );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(n2930), .D(n3017), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(n2928), .D(n3014), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n2930), .D(n3011), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(n2928), .D(n3008), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(n2929), .D(n3005), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(n2928), .D(n3002), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(n2929), .D(n2999), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(n2929), .D(n2996), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(n2929), .D(n2993), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(n2930), .D(n2990), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(n2927), .D(n3085), .Q(
        \REGISTERS[21][31] ) );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(n2925), .D(n3079), .Q(
        \REGISTERS[21][30] ) );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(n2927), .D(n3076), .Q(
        \REGISTERS[21][29] ) );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(n2925), .D(n3073), .Q(
        \REGISTERS[21][28] ) );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(n2927), .D(n3070), .Q(
        \REGISTERS[21][27] ) );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(n2925), .D(n3067), .Q(
        \REGISTERS[21][26] ) );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(n2925), .D(n3064), .Q(
        \REGISTERS[21][25] ) );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(n2925), .D(n3061), .Q(
        \REGISTERS[21][24] ) );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n2927), .D(n3058), .Q(
        \REGISTERS[21][23] ) );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n2925), .D(n3055), .Q(
        \REGISTERS[21][22] ) );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(n2925), .D(n3052), .Q(
        \REGISTERS[21][21] ) );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(n2926), .D(n3049), .Q(
        \REGISTERS[21][20] ) );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n2927), .D(n3046), .Q(
        \REGISTERS[21][19] ) );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(n2926), .D(n3043), .Q(
        \REGISTERS[21][18] ) );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n2926), .D(n3040), .Q(
        \REGISTERS[21][17] ) );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(n2926), .D(n3037), .Q(
        \REGISTERS[21][16] ) );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(n2925), .D(n3034), .Q(
        \REGISTERS[21][15] ) );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(n2926), .D(n3031), .Q(
        \REGISTERS[21][14] ) );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(n2926), .D(n3028), .Q(
        \REGISTERS[21][13] ) );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(n2926), .D(n3025), .Q(
        \REGISTERS[21][12] ) );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(n2927), .D(n3022), .Q(
        \REGISTERS[21][11] ) );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n2927), .D(n3019), .Q(
        \REGISTERS[21][10] ) );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(n2927), .D(n3016), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(n2925), .D(n3013), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n2927), .D(n3010), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(n2925), .D(n3007), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(n2926), .D(n3004), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(n2925), .D(n3001), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(n2926), .D(n2998), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(n2926), .D(n2995), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(n2926), .D(n2992), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(n2927), .D(n2989), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(n2924), .D(n3084), .Q(
        \REGISTERS[22][31] ) );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(n2922), .D(n3078), .Q(
        \REGISTERS[22][30] ) );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(n2924), .D(n3075), .Q(
        \REGISTERS[22][29] ) );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(n2922), .D(n3072), .Q(
        \REGISTERS[22][28] ) );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(n2924), .D(n3069), .Q(
        \REGISTERS[22][27] ) );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(n2922), .D(n3066), .Q(
        \REGISTERS[22][26] ) );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(n2922), .D(n3063), .Q(
        \REGISTERS[22][25] ) );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(n2922), .D(n3060), .Q(
        \REGISTERS[22][24] ) );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n2924), .D(n3057), .Q(
        \REGISTERS[22][23] ) );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n2922), .D(n3054), .Q(
        \REGISTERS[22][22] ) );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(n2922), .D(n3051), .Q(
        \REGISTERS[22][21] ) );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(n2923), .D(n3048), .Q(
        \REGISTERS[22][20] ) );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n2924), .D(n3045), .Q(
        \REGISTERS[22][19] ) );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(n2923), .D(n3042), .Q(
        \REGISTERS[22][18] ) );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n2923), .D(n3039), .Q(
        \REGISTERS[22][17] ) );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(n2923), .D(n3036), .Q(
        \REGISTERS[22][16] ) );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(n2922), .D(n3033), .Q(
        \REGISTERS[22][15] ) );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(n2923), .D(n3030), .Q(
        \REGISTERS[22][14] ) );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(n2923), .D(n3027), .Q(
        \REGISTERS[22][13] ) );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(n2923), .D(n3024), .Q(
        \REGISTERS[22][12] ) );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(n2924), .D(n3021), .Q(
        \REGISTERS[22][11] ) );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n2924), .D(n3018), .Q(
        \REGISTERS[22][10] ) );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(n2924), .D(n3015), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(n2922), .D(n3012), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n2924), .D(n3009), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(n2922), .D(n3006), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(n2923), .D(n3003), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(n2922), .D(n3000), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(n2923), .D(n2997), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(n2923), .D(n2994), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(n2923), .D(n2991), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(n2924), .D(n2988), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(n2921), .D(n3084), .Q(
        \REGISTERS[23][31] ) );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(n2919), .D(n3078), .Q(
        \REGISTERS[23][30] ) );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(n2921), .D(n3075), .Q(
        \REGISTERS[23][29] ) );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(n2919), .D(n3072), .Q(
        \REGISTERS[23][28] ) );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(n2921), .D(n3069), .Q(
        \REGISTERS[23][27] ) );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(n2919), .D(n3066), .Q(
        \REGISTERS[23][26] ) );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(n2919), .D(n3063), .Q(
        \REGISTERS[23][25] ) );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(n2919), .D(n3060), .Q(
        \REGISTERS[23][24] ) );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n2921), .D(n3057), .Q(
        \REGISTERS[23][23] ) );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n2919), .D(n3054), .Q(
        \REGISTERS[23][22] ) );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(n2919), .D(n3051), .Q(
        \REGISTERS[23][21] ) );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(n2920), .D(n3048), .Q(
        \REGISTERS[23][20] ) );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n2921), .D(n3045), .Q(
        \REGISTERS[23][19] ) );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(n2920), .D(n3042), .Q(
        \REGISTERS[23][18] ) );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n2920), .D(n3039), .Q(
        \REGISTERS[23][17] ) );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(n2920), .D(n3036), .Q(
        \REGISTERS[23][16] ) );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(n2919), .D(n3033), .Q(
        \REGISTERS[23][15] ) );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(n2920), .D(n3030), .Q(
        \REGISTERS[23][14] ) );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(n2920), .D(n3027), .Q(
        \REGISTERS[23][13] ) );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(n2920), .D(n3024), .Q(
        \REGISTERS[23][12] ) );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(n2921), .D(n3021), .Q(
        \REGISTERS[23][11] ) );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n2921), .D(n3018), .Q(
        \REGISTERS[23][10] ) );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(n2921), .D(n3015), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(n2919), .D(n3012), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n2921), .D(n3009), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(n2919), .D(n3006), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(n2920), .D(n3003), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(n2919), .D(n3000), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(n2920), .D(n2997), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(n2920), .D(n2994), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(n2920), .D(n2991), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(n2921), .D(n2988), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(n2918), .D(n3084), .Q(
        \REGISTERS[24][31] ) );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(n2916), .D(n3078), .Q(
        \REGISTERS[24][30] ) );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(n2918), .D(n3075), .Q(
        \REGISTERS[24][29] ) );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(n2916), .D(n3072), .Q(
        \REGISTERS[24][28] ) );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(n2918), .D(n3069), .Q(
        \REGISTERS[24][27] ) );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(n2916), .D(n3066), .Q(
        \REGISTERS[24][26] ) );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(n2916), .D(n3063), .Q(
        \REGISTERS[24][25] ) );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n2916), .D(n3060), .Q(
        \REGISTERS[24][24] ) );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n2918), .D(n3057), .Q(
        \REGISTERS[24][23] ) );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(n2916), .D(n3054), .Q(
        \REGISTERS[24][22] ) );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n2916), .D(n3051), .Q(
        \REGISTERS[24][21] ) );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n2917), .D(n3048), .Q(
        \REGISTERS[24][20] ) );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(n2918), .D(n3045), .Q(
        \REGISTERS[24][19] ) );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(n2917), .D(n3042), .Q(
        \REGISTERS[24][18] ) );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(n2917), .D(n3039), .Q(
        \REGISTERS[24][17] ) );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(n2917), .D(n3036), .Q(
        \REGISTERS[24][16] ) );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n2916), .D(n3033), .Q(
        \REGISTERS[24][15] ) );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(n2917), .D(n3030), .Q(
        \REGISTERS[24][14] ) );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(n2917), .D(n3027), .Q(
        \REGISTERS[24][13] ) );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(n2917), .D(n3024), .Q(
        \REGISTERS[24][12] ) );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(n2918), .D(n3021), .Q(
        \REGISTERS[24][11] ) );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(n2918), .D(n3018), .Q(
        \REGISTERS[24][10] ) );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(n2918), .D(n3015), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(n2916), .D(n3012), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(n2918), .D(n3009), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n2916), .D(n3006), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(n2917), .D(n3003), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(n2916), .D(n3000), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(n2917), .D(n2997), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(n2917), .D(n2994), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(n2917), .D(n2991), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(n2918), .D(n2988), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(n2915), .D(n3084), .Q(
        \REGISTERS[25][31] ) );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(n2913), .D(n3078), .Q(
        \REGISTERS[25][30] ) );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(n2915), .D(n3075), .Q(
        \REGISTERS[25][29] ) );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(n2913), .D(n3072), .Q(
        \REGISTERS[25][28] ) );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(n2915), .D(n3069), .Q(
        \REGISTERS[25][27] ) );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(n2913), .D(n3066), .Q(
        \REGISTERS[25][26] ) );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(n2913), .D(n3063), .Q(
        \REGISTERS[25][25] ) );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(n2913), .D(n3060), .Q(
        \REGISTERS[25][24] ) );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n2915), .D(n3057), .Q(
        \REGISTERS[25][23] ) );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n2913), .D(n3054), .Q(
        \REGISTERS[25][22] ) );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(n2913), .D(n3051), .Q(
        \REGISTERS[25][21] ) );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(n2914), .D(n3048), .Q(
        \REGISTERS[25][20] ) );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n2915), .D(n3045), .Q(
        \REGISTERS[25][19] ) );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(n2914), .D(n3042), .Q(
        \REGISTERS[25][18] ) );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n2914), .D(n3039), .Q(
        \REGISTERS[25][17] ) );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(n2914), .D(n3036), .Q(
        \REGISTERS[25][16] ) );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(n2913), .D(n3033), .Q(
        \REGISTERS[25][15] ) );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(n2914), .D(n3030), .Q(
        \REGISTERS[25][14] ) );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(n2914), .D(n3027), .Q(
        \REGISTERS[25][13] ) );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(n2914), .D(n3024), .Q(
        \REGISTERS[25][12] ) );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(n2915), .D(n3021), .Q(
        \REGISTERS[25][11] ) );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n2915), .D(n3018), .Q(
        \REGISTERS[25][10] ) );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(n2915), .D(n3015), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(n2913), .D(n3012), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n2915), .D(n3009), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(n2913), .D(n3006), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(n2914), .D(n3003), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(n2913), .D(n3000), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(n2914), .D(n2997), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(n2914), .D(n2994), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(n2914), .D(n2991), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(n2915), .D(n2988), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(n2912), .D(n3084), .Q(
        \REGISTERS[26][31] ) );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(n2910), .D(n3078), .Q(
        \REGISTERS[26][30] ) );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(n2912), .D(n3075), .Q(
        \REGISTERS[26][29] ) );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(n2910), .D(n3072), .Q(
        \REGISTERS[26][28] ) );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(n2912), .D(n3069), .Q(
        \REGISTERS[26][27] ) );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(n2910), .D(n3066), .Q(
        \REGISTERS[26][26] ) );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(n2910), .D(n3063), .Q(
        \REGISTERS[26][25] ) );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(n2910), .D(n3060), .Q(
        \REGISTERS[26][24] ) );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n2912), .D(n3057), .Q(
        \REGISTERS[26][23] ) );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n2910), .D(n3054), .Q(
        \REGISTERS[26][22] ) );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(n2910), .D(n3051), .Q(
        \REGISTERS[26][21] ) );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(n2911), .D(n3048), .Q(
        \REGISTERS[26][20] ) );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n2912), .D(n3045), .Q(
        \REGISTERS[26][19] ) );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(n2911), .D(n3042), .Q(
        \REGISTERS[26][18] ) );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n2911), .D(n3039), .Q(
        \REGISTERS[26][17] ) );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(n2911), .D(n3036), .Q(
        \REGISTERS[26][16] ) );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(n2910), .D(n3033), .Q(
        \REGISTERS[26][15] ) );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(n2911), .D(n3030), .Q(
        \REGISTERS[26][14] ) );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(n2911), .D(n3027), .Q(
        \REGISTERS[26][13] ) );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(n2911), .D(n3024), .Q(
        \REGISTERS[26][12] ) );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(n2912), .D(n3021), .Q(
        \REGISTERS[26][11] ) );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n2912), .D(n3018), .Q(
        \REGISTERS[26][10] ) );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(n2912), .D(n3015), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(n2910), .D(n3012), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n2912), .D(n3009), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(n2910), .D(n3006), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(n2911), .D(n3003), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(n2910), .D(n3000), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(n2911), .D(n2997), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(n2911), .D(n2994), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(n2911), .D(n2991), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(n2912), .D(n2988), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(n2909), .D(n3084), .Q(
        \REGISTERS[27][31] ) );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(n2907), .D(n3078), .Q(
        \REGISTERS[27][30] ) );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(n2909), .D(n3075), .Q(
        \REGISTERS[27][29] ) );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(n2907), .D(n3072), .Q(
        \REGISTERS[27][28] ) );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(n2909), .D(n3069), .Q(
        \REGISTERS[27][27] ) );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(n2907), .D(n3066), .Q(
        \REGISTERS[27][26] ) );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(n2907), .D(n3063), .Q(
        \REGISTERS[27][25] ) );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(n2907), .D(n3060), .Q(
        \REGISTERS[27][24] ) );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n2909), .D(n3057), .Q(
        \REGISTERS[27][23] ) );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n2907), .D(n3054), .Q(
        \REGISTERS[27][22] ) );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(n2907), .D(n3051), .Q(
        \REGISTERS[27][21] ) );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(n2908), .D(n3048), .Q(
        \REGISTERS[27][20] ) );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n2909), .D(n3045), .Q(
        \REGISTERS[27][19] ) );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(n2908), .D(n3042), .Q(
        \REGISTERS[27][18] ) );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n2908), .D(n3039), .Q(
        \REGISTERS[27][17] ) );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(n2908), .D(n3036), .Q(
        \REGISTERS[27][16] ) );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(n2907), .D(n3033), .Q(
        \REGISTERS[27][15] ) );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(n2908), .D(n3030), .Q(
        \REGISTERS[27][14] ) );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(n2908), .D(n3027), .Q(
        \REGISTERS[27][13] ) );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(n2908), .D(n3024), .Q(
        \REGISTERS[27][12] ) );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(n2909), .D(n3021), .Q(
        \REGISTERS[27][11] ) );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n2909), .D(n3018), .Q(
        \REGISTERS[27][10] ) );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(n2909), .D(n3015), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(n2907), .D(n3012), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n2909), .D(n3009), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(n2907), .D(n3006), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(n2908), .D(n3003), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(n2907), .D(n3000), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(n2908), .D(n2997), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(n2908), .D(n2994), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(n2908), .D(n2991), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(n2909), .D(n2988), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(n2906), .D(n3084), .Q(
        \REGISTERS[28][31] ) );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(n2904), .D(n3078), .Q(
        \REGISTERS[28][30] ) );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(n2906), .D(n3075), .Q(
        \REGISTERS[28][29] ) );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(n2904), .D(n3072), .Q(
        \REGISTERS[28][28] ) );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(n2906), .D(n3069), .Q(
        \REGISTERS[28][27] ) );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(n2904), .D(n3066), .Q(
        \REGISTERS[28][26] ) );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(n2904), .D(n3063), .Q(
        \REGISTERS[28][25] ) );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(n2904), .D(n3060), .Q(
        \REGISTERS[28][24] ) );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n2906), .D(n3057), .Q(
        \REGISTERS[28][23] ) );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n2904), .D(n3054), .Q(
        \REGISTERS[28][22] ) );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(n2904), .D(n3051), .Q(
        \REGISTERS[28][21] ) );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(n2905), .D(n3048), .Q(
        \REGISTERS[28][20] ) );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n2906), .D(n3045), .Q(
        \REGISTERS[28][19] ) );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(n2905), .D(n3042), .Q(
        \REGISTERS[28][18] ) );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n2905), .D(n3039), .Q(
        \REGISTERS[28][17] ) );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(n2905), .D(n3036), .Q(
        \REGISTERS[28][16] ) );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(n2904), .D(n3033), .Q(
        \REGISTERS[28][15] ) );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(n2905), .D(n3030), .Q(
        \REGISTERS[28][14] ) );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(n2905), .D(n3027), .Q(
        \REGISTERS[28][13] ) );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(n2905), .D(n3024), .Q(
        \REGISTERS[28][12] ) );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(n2906), .D(n3021), .Q(
        \REGISTERS[28][11] ) );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n2906), .D(n3018), .Q(
        \REGISTERS[28][10] ) );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(n2906), .D(n3015), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(n2904), .D(n3012), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n2906), .D(n3009), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(n2904), .D(n3006), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(n2905), .D(n3003), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(n2904), .D(n3000), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(n2905), .D(n2997), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(n2905), .D(n2994), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(n2905), .D(n2991), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(n2906), .D(n2988), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(n2903), .D(n3084), .Q(
        \REGISTERS[29][31] ) );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(n2901), .D(n3078), .Q(
        \REGISTERS[29][30] ) );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(n2903), .D(n3075), .Q(
        \REGISTERS[29][29] ) );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(n2901), .D(n3072), .Q(
        \REGISTERS[29][28] ) );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(n2903), .D(n3069), .Q(
        \REGISTERS[29][27] ) );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(n2901), .D(n3066), .Q(
        \REGISTERS[29][26] ) );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(n2901), .D(n3063), .Q(
        \REGISTERS[29][25] ) );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(n2901), .D(n3060), .Q(
        \REGISTERS[29][24] ) );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n2903), .D(n3057), .Q(
        \REGISTERS[29][23] ) );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n2901), .D(n3054), .Q(
        \REGISTERS[29][22] ) );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(n2901), .D(n3051), .Q(
        \REGISTERS[29][21] ) );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(n2902), .D(n3048), .Q(
        \REGISTERS[29][20] ) );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n2903), .D(n3045), .Q(
        \REGISTERS[29][19] ) );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(n2902), .D(n3042), .Q(
        \REGISTERS[29][18] ) );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n2902), .D(n3039), .Q(
        \REGISTERS[29][17] ) );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(n2902), .D(n3036), .Q(
        \REGISTERS[29][16] ) );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(n2901), .D(n3033), .Q(
        \REGISTERS[29][15] ) );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(n2902), .D(n3030), .Q(
        \REGISTERS[29][14] ) );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(n2902), .D(n3027), .Q(
        \REGISTERS[29][13] ) );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(n2902), .D(n3024), .Q(
        \REGISTERS[29][12] ) );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(n2903), .D(n3021), .Q(
        \REGISTERS[29][11] ) );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n2903), .D(n3018), .Q(
        \REGISTERS[29][10] ) );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(n2903), .D(n3015), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(n2901), .D(n3012), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n2903), .D(n3009), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(n2901), .D(n3006), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(n2902), .D(n3003), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(n2901), .D(n3000), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(n2902), .D(n2997), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(n2902), .D(n2994), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(n2902), .D(n2991), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(n2903), .D(n2988), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(n2900), .D(n3084), .Q(
        \REGISTERS[30][31] ) );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(n2898), .D(n3078), .Q(
        \REGISTERS[30][30] ) );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(n2900), .D(n3075), .Q(
        \REGISTERS[30][29] ) );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(n2898), .D(n3072), .Q(
        \REGISTERS[30][28] ) );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(n2900), .D(n3069), .Q(
        \REGISTERS[30][27] ) );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(n2898), .D(n3066), .Q(
        \REGISTERS[30][26] ) );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(n2898), .D(n3063), .Q(
        \REGISTERS[30][25] ) );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(n2898), .D(n3060), .Q(
        \REGISTERS[30][24] ) );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n2900), .D(n3057), .Q(
        \REGISTERS[30][23] ) );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n2898), .D(n3054), .Q(
        \REGISTERS[30][22] ) );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(n2898), .D(n3051), .Q(
        \REGISTERS[30][21] ) );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(n2899), .D(n3048), .Q(
        \REGISTERS[30][20] ) );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n2900), .D(n3045), .Q(
        \REGISTERS[30][19] ) );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(n2899), .D(n3042), .Q(
        \REGISTERS[30][18] ) );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n2899), .D(n3039), .Q(
        \REGISTERS[30][17] ) );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(n2899), .D(n3036), .Q(
        \REGISTERS[30][16] ) );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(n2898), .D(n3033), .Q(
        \REGISTERS[30][15] ) );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(n2899), .D(n3030), .Q(
        \REGISTERS[30][14] ) );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(n2899), .D(n3027), .Q(
        \REGISTERS[30][13] ) );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(n2899), .D(n3024), .Q(
        \REGISTERS[30][12] ) );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(n2900), .D(n3021), .Q(
        \REGISTERS[30][11] ) );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n2900), .D(n3018), .Q(
        \REGISTERS[30][10] ) );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(n2900), .D(n3015), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(n2898), .D(n3012), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n2900), .D(n3009), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(n2898), .D(n3006), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(n2899), .D(n3003), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(n2898), .D(n3000), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(n2899), .D(n2997), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(n2899), .D(n2994), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(n2899), .D(n2991), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(n2900), .D(n2988), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(n2897), .D(n3084), .Q(
        \REGISTERS[31][31] ) );
  DLH_X1 \OUT2_reg[31]  ( .G(n3091), .D(N4529), .Q(OUT2[31]) );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(n2895), .D(n3078), .Q(
        \REGISTERS[31][30] ) );
  DLH_X1 \OUT2_reg[30]  ( .G(n3091), .D(N4527), .Q(OUT2[30]) );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(n2897), .D(n3075), .Q(
        \REGISTERS[31][29] ) );
  DLH_X1 \OUT2_reg[29]  ( .G(n3091), .D(N4525), .Q(OUT2[29]) );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(n2895), .D(n3072), .Q(
        \REGISTERS[31][28] ) );
  DLH_X1 \OUT2_reg[28]  ( .G(n3092), .D(N4523), .Q(OUT2[28]) );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(n2897), .D(n3069), .Q(
        \REGISTERS[31][27] ) );
  DLH_X1 \OUT2_reg[27]  ( .G(n3091), .D(N4521), .Q(OUT2[27]) );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(n2895), .D(n3066), .Q(
        \REGISTERS[31][26] ) );
  DLH_X1 \OUT2_reg[26]  ( .G(n3092), .D(N4519), .Q(OUT2[26]) );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(n2895), .D(n3063), .Q(
        \REGISTERS[31][25] ) );
  DLH_X1 \OUT2_reg[25]  ( .G(n3092), .D(N4517), .Q(OUT2[25]) );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(n2895), .D(n3060), .Q(
        \REGISTERS[31][24] ) );
  DLH_X1 \OUT2_reg[24]  ( .G(n3092), .D(N4515), .Q(OUT2[24]) );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(n2897), .D(n3057), .Q(
        \REGISTERS[31][23] ) );
  DLH_X1 \OUT2_reg[23]  ( .G(n3091), .D(N4513), .Q(OUT2[23]) );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(n2895), .D(n3054), .Q(
        \REGISTERS[31][22] ) );
  DLH_X1 \OUT2_reg[22]  ( .G(n3091), .D(N4511), .Q(OUT2[22]) );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n2895), .D(n3051), .Q(
        \REGISTERS[31][21] ) );
  DLH_X1 \OUT2_reg[21]  ( .G(n3092), .D(N4509), .Q(OUT2[21]) );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(n2896), .D(n3048), .Q(
        \REGISTERS[31][20] ) );
  DLH_X1 \OUT2_reg[20]  ( .G(n3092), .D(N4507), .Q(OUT2[20]) );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n2897), .D(n3045), .Q(
        \REGISTERS[31][19] ) );
  DLH_X1 \OUT2_reg[19]  ( .G(n3091), .D(N4505), .Q(OUT2[19]) );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(n2896), .D(n3042), .Q(
        \REGISTERS[31][18] ) );
  DLH_X1 \OUT2_reg[18]  ( .G(n3090), .D(N4503), .Q(OUT2[18]) );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n2896), .D(n3039), .Q(
        \REGISTERS[31][17] ) );
  DLH_X1 \OUT2_reg[17]  ( .G(n3090), .D(N4501), .Q(OUT2[17]) );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(n2896), .D(n3036), .Q(
        \REGISTERS[31][16] ) );
  DLH_X1 \OUT2_reg[16]  ( .G(n3090), .D(N4499), .Q(OUT2[16]) );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(n2895), .D(n3033), .Q(
        \REGISTERS[31][15] ) );
  DLH_X1 \OUT2_reg[15]  ( .G(n3092), .D(N4497), .Q(OUT2[15]) );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(n2896), .D(n3030), .Q(
        \REGISTERS[31][14] ) );
  DLH_X1 \OUT2_reg[14]  ( .G(n3090), .D(N4495), .Q(OUT2[14]) );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(n2896), .D(n3027), .Q(
        \REGISTERS[31][13] ) );
  DLH_X1 \OUT2_reg[13]  ( .G(n3090), .D(N4493), .Q(OUT2[13]) );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(n2896), .D(n3024), .Q(
        \REGISTERS[31][12] ) );
  DLH_X1 \OUT2_reg[12]  ( .G(n3090), .D(N4491), .Q(OUT2[12]) );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n2897), .D(n3021), .Q(
        \REGISTERS[31][11] ) );
  DLH_X1 \OUT2_reg[11]  ( .G(n3091), .D(N4489), .Q(OUT2[11]) );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n2897), .D(n3018), .Q(
        \REGISTERS[31][10] ) );
  DLH_X1 \OUT2_reg[10]  ( .G(n3091), .D(N4487), .Q(OUT2[10]) );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(n2897), .D(n3015), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \OUT2_reg[9]  ( .G(n3091), .D(N4485), .Q(OUT2[9]) );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(n2895), .D(n3012), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \OUT2_reg[8]  ( .G(n3092), .D(N4483), .Q(OUT2[8]) );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(n2897), .D(n3009), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \OUT2_reg[7]  ( .G(n3091), .D(N4481), .Q(OUT2[7]) );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(n2895), .D(n3006), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \OUT2_reg[6]  ( .G(n3092), .D(N4479), .Q(OUT2[6]) );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(n2896), .D(n3003), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \OUT2_reg[5]  ( .G(n3090), .D(N4477), .Q(OUT2[5]) );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(n2895), .D(n3000), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \OUT2_reg[4]  ( .G(n3092), .D(N4475), .Q(OUT2[4]) );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(n2896), .D(n2997), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \OUT2_reg[3]  ( .G(n3090), .D(N4473), .Q(OUT2[3]) );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(n2896), .D(n2994), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \OUT2_reg[2]  ( .G(n3090), .D(N4471), .Q(OUT2[2]) );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(n2896), .D(n2991), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \OUT2_reg[1]  ( .G(n3090), .D(N4469), .Q(OUT2[1]) );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n2897), .D(n2988), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUT2_reg[0]  ( .G(n3090), .D(N4467), .Q(OUT2[0]) );
  DLH_X1 \OUT1_reg[31]  ( .G(n3088), .D(N4465), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n3088), .D(N4463), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n3088), .D(N4461), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n3089), .D(N4459), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n3088), .D(N4457), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n3089), .D(N4455), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n3089), .D(N4453), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n3089), .D(N4451), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n3088), .D(N4449), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n3089), .D(N4447), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n3089), .D(N4445), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n3088), .D(N4443), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n3088), .D(N4441), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n3087), .D(N4439), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n3087), .D(N4437), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n3087), .D(N4435), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n3089), .D(N4433), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n3087), .D(N4431), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n3087), .D(N4429), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n3087), .D(N4427), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n3088), .D(N4425), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n3088), .D(N4423), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n3088), .D(N4421), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n3089), .D(N4419), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n3088), .D(N4417), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n3089), .D(N4415), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n3087), .D(N4413), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n3089), .D(N4411), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n3087), .D(N4409), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n3087), .D(N4407), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n3087), .D(N4405), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n3087), .D(N4403), .Q(OUT1[0]) );
  NAND3_X1 U1901 ( .A1(ADD_WR[3]), .A2(n535), .A3(ADD_WR[4]), .ZN(n526) );
  NAND3_X1 U1902 ( .A1(n535), .A2(n537), .A3(ADD_WR[4]), .ZN(n536) );
  NAND3_X1 U1903 ( .A1(n535), .A2(n539), .A3(ADD_WR[3]), .ZN(n538) );
  NAND3_X1 U1904 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n527)
         );
  NAND3_X1 U1905 ( .A1(ADD_WR[1]), .A2(n541), .A3(ADD_WR[2]), .ZN(n528) );
  NAND3_X1 U1906 ( .A1(ADD_WR[0]), .A2(n542), .A3(ADD_WR[2]), .ZN(n529) );
  NAND3_X1 U1907 ( .A1(n541), .A2(n542), .A3(ADD_WR[2]), .ZN(n530) );
  NAND3_X1 U1908 ( .A1(ADD_WR[0]), .A2(n543), .A3(ADD_WR[1]), .ZN(n531) );
  NAND3_X1 U1909 ( .A1(n541), .A2(n543), .A3(ADD_WR[1]), .ZN(n532) );
  NAND3_X1 U1910 ( .A1(n542), .A2(n543), .A3(ADD_WR[0]), .ZN(n533) );
  NAND3_X1 U1911 ( .A1(n537), .A2(n539), .A3(n535), .ZN(n540) );
  NAND3_X1 U1912 ( .A1(n542), .A2(n543), .A3(n541), .ZN(n534) );
  BUF_X1 U3 ( .A(n2509), .Z(n3082) );
  BUF_X1 U4 ( .A(n2509), .Z(n3081) );
  BUF_X1 U5 ( .A(n2509), .Z(n3083) );
  OAI21_X1 U6 ( .B1(n534), .B2(n540), .A(n3095), .ZN(n2509) );
  BUF_X1 U7 ( .A(n557), .Z(n2886) );
  BUF_X1 U8 ( .A(n564), .Z(n2874) );
  BUF_X1 U9 ( .A(n571), .Z(n2862) );
  BUF_X1 U10 ( .A(n578), .Z(n2850) );
  BUF_X1 U11 ( .A(n589), .Z(n2838) );
  BUF_X1 U12 ( .A(n596), .Z(n2826) );
  BUF_X1 U13 ( .A(n603), .Z(n2814) );
  BUF_X1 U14 ( .A(n610), .Z(n2802) );
  BUF_X1 U15 ( .A(n557), .Z(n2887) );
  BUF_X1 U16 ( .A(n564), .Z(n2875) );
  BUF_X1 U17 ( .A(n571), .Z(n2863) );
  BUF_X1 U18 ( .A(n578), .Z(n2851) );
  BUF_X1 U19 ( .A(n589), .Z(n2839) );
  BUF_X1 U20 ( .A(n596), .Z(n2827) );
  BUF_X1 U21 ( .A(n603), .Z(n2815) );
  BUF_X1 U22 ( .A(n610), .Z(n2803) );
  BUF_X1 U23 ( .A(n552), .Z(n2892) );
  BUF_X1 U24 ( .A(n559), .Z(n2880) );
  BUF_X1 U25 ( .A(n566), .Z(n2868) );
  BUF_X1 U26 ( .A(n573), .Z(n2856) );
  BUF_X1 U27 ( .A(n584), .Z(n2844) );
  BUF_X1 U28 ( .A(n591), .Z(n2832) );
  BUF_X1 U29 ( .A(n598), .Z(n2820) );
  BUF_X1 U30 ( .A(n605), .Z(n2808) );
  BUF_X1 U31 ( .A(n552), .Z(n2893) );
  BUF_X1 U32 ( .A(n559), .Z(n2881) );
  BUF_X1 U33 ( .A(n566), .Z(n2869) );
  BUF_X1 U34 ( .A(n573), .Z(n2857) );
  BUF_X1 U35 ( .A(n584), .Z(n2845) );
  BUF_X1 U36 ( .A(n591), .Z(n2833) );
  BUF_X1 U37 ( .A(n598), .Z(n2821) );
  BUF_X1 U38 ( .A(n605), .Z(n2809) );
  BUF_X1 U39 ( .A(n558), .Z(n2883) );
  BUF_X1 U40 ( .A(n565), .Z(n2871) );
  BUF_X1 U41 ( .A(n572), .Z(n2859) );
  BUF_X1 U42 ( .A(n579), .Z(n2847) );
  BUF_X1 U43 ( .A(n590), .Z(n2835) );
  BUF_X1 U44 ( .A(n597), .Z(n2823) );
  BUF_X1 U45 ( .A(n604), .Z(n2811) );
  BUF_X1 U46 ( .A(n611), .Z(n2799) );
  BUF_X1 U47 ( .A(n558), .Z(n2884) );
  BUF_X1 U48 ( .A(n565), .Z(n2872) );
  BUF_X1 U49 ( .A(n572), .Z(n2860) );
  BUF_X1 U50 ( .A(n579), .Z(n2848) );
  BUF_X1 U51 ( .A(n590), .Z(n2836) );
  BUF_X1 U52 ( .A(n597), .Z(n2824) );
  BUF_X1 U53 ( .A(n604), .Z(n2812) );
  BUF_X1 U54 ( .A(n611), .Z(n2800) );
  BUF_X1 U55 ( .A(n1689), .Z(n2793) );
  BUF_X1 U56 ( .A(n1694), .Z(n2781) );
  BUF_X1 U57 ( .A(n1699), .Z(n2769) );
  BUF_X1 U58 ( .A(n1704), .Z(n2757) );
  BUF_X1 U59 ( .A(n1713), .Z(n2745) );
  BUF_X1 U60 ( .A(n1718), .Z(n2733) );
  BUF_X1 U61 ( .A(n1723), .Z(n2721) );
  BUF_X1 U62 ( .A(n1728), .Z(n2709) );
  BUF_X1 U63 ( .A(n1689), .Z(n2794) );
  BUF_X1 U64 ( .A(n1694), .Z(n2782) );
  BUF_X1 U65 ( .A(n1699), .Z(n2770) );
  BUF_X1 U66 ( .A(n1704), .Z(n2758) );
  BUF_X1 U67 ( .A(n1713), .Z(n2746) );
  BUF_X1 U68 ( .A(n1718), .Z(n2734) );
  BUF_X1 U69 ( .A(n1723), .Z(n2722) );
  BUF_X1 U70 ( .A(n1728), .Z(n2710) );
  BUF_X1 U71 ( .A(n1691), .Z(n2790) );
  BUF_X1 U72 ( .A(n1696), .Z(n2778) );
  BUF_X1 U73 ( .A(n1701), .Z(n2766) );
  BUF_X1 U74 ( .A(n1706), .Z(n2754) );
  BUF_X1 U75 ( .A(n1715), .Z(n2742) );
  BUF_X1 U76 ( .A(n1720), .Z(n2730) );
  BUF_X1 U77 ( .A(n1725), .Z(n2718) );
  BUF_X1 U78 ( .A(n1730), .Z(n2706) );
  BUF_X1 U79 ( .A(n1691), .Z(n2791) );
  BUF_X1 U80 ( .A(n1696), .Z(n2779) );
  BUF_X1 U81 ( .A(n1701), .Z(n2767) );
  BUF_X1 U82 ( .A(n1706), .Z(n2755) );
  BUF_X1 U83 ( .A(n1715), .Z(n2743) );
  BUF_X1 U84 ( .A(n1720), .Z(n2731) );
  BUF_X1 U85 ( .A(n1725), .Z(n2719) );
  BUF_X1 U86 ( .A(n1730), .Z(n2707) );
  BUF_X1 U87 ( .A(n1688), .Z(n2796) );
  BUF_X1 U88 ( .A(n1693), .Z(n2784) );
  BUF_X1 U89 ( .A(n1698), .Z(n2772) );
  BUF_X1 U90 ( .A(n1703), .Z(n2760) );
  BUF_X1 U91 ( .A(n1712), .Z(n2748) );
  BUF_X1 U92 ( .A(n1717), .Z(n2736) );
  BUF_X1 U93 ( .A(n1722), .Z(n2724) );
  BUF_X1 U94 ( .A(n1727), .Z(n2712) );
  BUF_X1 U95 ( .A(n1688), .Z(n2797) );
  BUF_X1 U96 ( .A(n1693), .Z(n2785) );
  BUF_X1 U97 ( .A(n1698), .Z(n2773) );
  BUF_X1 U98 ( .A(n1703), .Z(n2761) );
  BUF_X1 U99 ( .A(n1712), .Z(n2749) );
  BUF_X1 U100 ( .A(n1717), .Z(n2737) );
  BUF_X1 U101 ( .A(n1722), .Z(n2725) );
  BUF_X1 U102 ( .A(n1727), .Z(n2713) );
  BUF_X1 U103 ( .A(n557), .Z(n2888) );
  BUF_X1 U104 ( .A(n564), .Z(n2876) );
  BUF_X1 U105 ( .A(n578), .Z(n2852) );
  BUF_X1 U106 ( .A(n589), .Z(n2840) );
  BUF_X1 U107 ( .A(n603), .Z(n2816) );
  BUF_X1 U108 ( .A(n610), .Z(n2804) );
  BUF_X1 U109 ( .A(n552), .Z(n2894) );
  BUF_X1 U110 ( .A(n559), .Z(n2882) );
  BUF_X1 U111 ( .A(n571), .Z(n2864) );
  BUF_X1 U112 ( .A(n596), .Z(n2828) );
  BUF_X1 U113 ( .A(n566), .Z(n2870) );
  BUF_X1 U114 ( .A(n573), .Z(n2858) );
  BUF_X1 U115 ( .A(n584), .Z(n2846) );
  BUF_X1 U116 ( .A(n591), .Z(n2834) );
  BUF_X1 U117 ( .A(n598), .Z(n2822) );
  BUF_X1 U118 ( .A(n605), .Z(n2810) );
  BUF_X1 U119 ( .A(n558), .Z(n2885) );
  BUF_X1 U120 ( .A(n565), .Z(n2873) );
  BUF_X1 U121 ( .A(n572), .Z(n2861) );
  BUF_X1 U122 ( .A(n579), .Z(n2849) );
  BUF_X1 U123 ( .A(n590), .Z(n2837) );
  BUF_X1 U124 ( .A(n597), .Z(n2825) );
  BUF_X1 U125 ( .A(n604), .Z(n2813) );
  BUF_X1 U126 ( .A(n611), .Z(n2801) );
  BUF_X1 U127 ( .A(n554), .Z(n2889) );
  BUF_X1 U128 ( .A(n561), .Z(n2877) );
  BUF_X1 U129 ( .A(n568), .Z(n2865) );
  BUF_X1 U130 ( .A(n575), .Z(n2853) );
  BUF_X1 U131 ( .A(n586), .Z(n2841) );
  BUF_X1 U132 ( .A(n593), .Z(n2829) );
  BUF_X1 U133 ( .A(n600), .Z(n2817) );
  BUF_X1 U134 ( .A(n607), .Z(n2805) );
  BUF_X1 U135 ( .A(n554), .Z(n2890) );
  BUF_X1 U136 ( .A(n561), .Z(n2878) );
  BUF_X1 U137 ( .A(n568), .Z(n2866) );
  BUF_X1 U138 ( .A(n575), .Z(n2854) );
  BUF_X1 U139 ( .A(n586), .Z(n2842) );
  BUF_X1 U140 ( .A(n593), .Z(n2830) );
  BUF_X1 U141 ( .A(n600), .Z(n2818) );
  BUF_X1 U142 ( .A(n607), .Z(n2806) );
  BUF_X1 U143 ( .A(n1692), .Z(n2788) );
  BUF_X1 U144 ( .A(n1697), .Z(n2776) );
  BUF_X1 U145 ( .A(n1702), .Z(n2764) );
  BUF_X1 U146 ( .A(n1707), .Z(n2752) );
  BUF_X1 U147 ( .A(n1716), .Z(n2740) );
  BUF_X1 U148 ( .A(n1721), .Z(n2728) );
  BUF_X1 U149 ( .A(n1726), .Z(n2716) );
  BUF_X1 U150 ( .A(n1731), .Z(n2704) );
  BUF_X1 U151 ( .A(n1692), .Z(n2787) );
  BUF_X1 U152 ( .A(n1697), .Z(n2775) );
  BUF_X1 U153 ( .A(n1702), .Z(n2763) );
  BUF_X1 U154 ( .A(n1707), .Z(n2751) );
  BUF_X1 U155 ( .A(n1716), .Z(n2739) );
  BUF_X1 U156 ( .A(n1721), .Z(n2727) );
  BUF_X1 U157 ( .A(n1726), .Z(n2715) );
  BUF_X1 U158 ( .A(n1731), .Z(n2703) );
  BUF_X1 U159 ( .A(n1713), .Z(n2747) );
  BUF_X1 U160 ( .A(n1718), .Z(n2735) );
  BUF_X1 U161 ( .A(n1723), .Z(n2723) );
  BUF_X1 U162 ( .A(n1728), .Z(n2711) );
  BUF_X1 U163 ( .A(n1689), .Z(n2795) );
  BUF_X1 U164 ( .A(n1694), .Z(n2783) );
  BUF_X1 U165 ( .A(n1699), .Z(n2771) );
  BUF_X1 U166 ( .A(n1704), .Z(n2759) );
  BUF_X1 U167 ( .A(n1691), .Z(n2792) );
  BUF_X1 U168 ( .A(n1696), .Z(n2780) );
  BUF_X1 U169 ( .A(n1701), .Z(n2768) );
  BUF_X1 U170 ( .A(n1706), .Z(n2756) );
  BUF_X1 U171 ( .A(n1715), .Z(n2744) );
  BUF_X1 U172 ( .A(n1720), .Z(n2732) );
  BUF_X1 U173 ( .A(n1725), .Z(n2720) );
  BUF_X1 U174 ( .A(n1730), .Z(n2708) );
  BUF_X1 U175 ( .A(n1712), .Z(n2750) );
  BUF_X1 U176 ( .A(n1717), .Z(n2738) );
  BUF_X1 U177 ( .A(n1722), .Z(n2726) );
  BUF_X1 U178 ( .A(n1727), .Z(n2714) );
  BUF_X1 U179 ( .A(n1688), .Z(n2798) );
  BUF_X1 U180 ( .A(n1693), .Z(n2786) );
  BUF_X1 U181 ( .A(n1698), .Z(n2774) );
  BUF_X1 U182 ( .A(n1703), .Z(n2762) );
  BUF_X1 U183 ( .A(n554), .Z(n2891) );
  BUF_X1 U184 ( .A(n561), .Z(n2879) );
  BUF_X1 U185 ( .A(n568), .Z(n2867) );
  BUF_X1 U186 ( .A(n575), .Z(n2855) );
  BUF_X1 U187 ( .A(n586), .Z(n2843) );
  BUF_X1 U188 ( .A(n593), .Z(n2831) );
  BUF_X1 U189 ( .A(n600), .Z(n2819) );
  BUF_X1 U190 ( .A(n607), .Z(n2807) );
  BUF_X1 U191 ( .A(n1692), .Z(n2789) );
  BUF_X1 U192 ( .A(n1697), .Z(n2777) );
  BUF_X1 U193 ( .A(n1702), .Z(n2765) );
  BUF_X1 U194 ( .A(n1707), .Z(n2753) );
  BUF_X1 U195 ( .A(n1716), .Z(n2741) );
  BUF_X1 U196 ( .A(n1721), .Z(n2729) );
  BUF_X1 U197 ( .A(n1726), .Z(n2717) );
  BUF_X1 U198 ( .A(n1731), .Z(n2705) );
  BUF_X1 U199 ( .A(n2695), .Z(n2896) );
  BUF_X1 U200 ( .A(n2695), .Z(n2895) );
  BUF_X1 U201 ( .A(n2692), .Z(n2899) );
  BUF_X1 U202 ( .A(n2692), .Z(n2898) );
  BUF_X1 U203 ( .A(n2689), .Z(n2902) );
  BUF_X1 U204 ( .A(n2689), .Z(n2901) );
  BUF_X1 U205 ( .A(n2686), .Z(n2905) );
  BUF_X1 U206 ( .A(n2686), .Z(n2904) );
  BUF_X1 U207 ( .A(n2683), .Z(n2908) );
  BUF_X1 U208 ( .A(n2683), .Z(n2907) );
  BUF_X1 U209 ( .A(n2680), .Z(n2911) );
  BUF_X1 U210 ( .A(n2680), .Z(n2910) );
  BUF_X1 U211 ( .A(n2677), .Z(n2914) );
  BUF_X1 U212 ( .A(n2677), .Z(n2913) );
  BUF_X1 U213 ( .A(n2674), .Z(n2917) );
  BUF_X1 U214 ( .A(n2674), .Z(n2916) );
  BUF_X1 U215 ( .A(n2671), .Z(n2920) );
  BUF_X1 U216 ( .A(n2671), .Z(n2919) );
  BUF_X1 U217 ( .A(n2668), .Z(n2923) );
  BUF_X1 U218 ( .A(n2668), .Z(n2922) );
  BUF_X1 U219 ( .A(n2665), .Z(n2926) );
  BUF_X1 U220 ( .A(n2665), .Z(n2925) );
  BUF_X1 U221 ( .A(n2662), .Z(n2929) );
  BUF_X1 U222 ( .A(n2662), .Z(n2928) );
  BUF_X1 U223 ( .A(n2659), .Z(n2932) );
  BUF_X1 U224 ( .A(n2659), .Z(n2931) );
  BUF_X1 U225 ( .A(n2656), .Z(n2935) );
  BUF_X1 U226 ( .A(n2656), .Z(n2934) );
  BUF_X1 U227 ( .A(n2653), .Z(n2938) );
  BUF_X1 U228 ( .A(n2653), .Z(n2937) );
  BUF_X1 U229 ( .A(n2650), .Z(n2941) );
  BUF_X1 U230 ( .A(n2650), .Z(n2940) );
  BUF_X1 U231 ( .A(n2647), .Z(n2944) );
  BUF_X1 U232 ( .A(n2647), .Z(n2943) );
  BUF_X1 U233 ( .A(n2644), .Z(n2947) );
  BUF_X1 U234 ( .A(n2644), .Z(n2946) );
  BUF_X1 U235 ( .A(n2641), .Z(n2950) );
  BUF_X1 U236 ( .A(n2641), .Z(n2949) );
  BUF_X1 U237 ( .A(n2638), .Z(n2953) );
  BUF_X1 U238 ( .A(n2638), .Z(n2952) );
  BUF_X1 U239 ( .A(n2635), .Z(n2956) );
  BUF_X1 U240 ( .A(n2635), .Z(n2955) );
  BUF_X1 U241 ( .A(n2632), .Z(n2959) );
  BUF_X1 U242 ( .A(n2632), .Z(n2958) );
  BUF_X1 U243 ( .A(n2629), .Z(n2962) );
  BUF_X1 U244 ( .A(n2629), .Z(n2961) );
  BUF_X1 U245 ( .A(n2626), .Z(n2965) );
  BUF_X1 U246 ( .A(n2626), .Z(n2964) );
  BUF_X1 U247 ( .A(n2623), .Z(n2968) );
  BUF_X1 U248 ( .A(n2623), .Z(n2967) );
  BUF_X1 U249 ( .A(n2620), .Z(n2971) );
  BUF_X1 U250 ( .A(n2620), .Z(n2970) );
  BUF_X1 U251 ( .A(n2617), .Z(n2974) );
  BUF_X1 U252 ( .A(n2617), .Z(n2973) );
  BUF_X1 U253 ( .A(n2614), .Z(n2977) );
  BUF_X1 U254 ( .A(n2614), .Z(n2976) );
  BUF_X1 U255 ( .A(n2611), .Z(n2980) );
  BUF_X1 U256 ( .A(n2611), .Z(n2979) );
  BUF_X1 U257 ( .A(n2608), .Z(n2983) );
  BUF_X1 U258 ( .A(n2608), .Z(n2982) );
  BUF_X1 U259 ( .A(n2605), .Z(n2986) );
  BUF_X1 U260 ( .A(n2605), .Z(n2985) );
  BUF_X1 U261 ( .A(n2695), .Z(n2897) );
  BUF_X1 U262 ( .A(n2692), .Z(n2900) );
  BUF_X1 U263 ( .A(n2689), .Z(n2903) );
  BUF_X1 U264 ( .A(n2686), .Z(n2906) );
  BUF_X1 U265 ( .A(n2683), .Z(n2909) );
  BUF_X1 U266 ( .A(n2680), .Z(n2912) );
  BUF_X1 U267 ( .A(n2677), .Z(n2915) );
  BUF_X1 U268 ( .A(n2674), .Z(n2918) );
  BUF_X1 U269 ( .A(n2671), .Z(n2921) );
  BUF_X1 U270 ( .A(n2668), .Z(n2924) );
  BUF_X1 U271 ( .A(n2665), .Z(n2927) );
  BUF_X1 U272 ( .A(n2662), .Z(n2930) );
  BUF_X1 U273 ( .A(n2659), .Z(n2933) );
  BUF_X1 U274 ( .A(n2656), .Z(n2936) );
  BUF_X1 U275 ( .A(n2653), .Z(n2939) );
  BUF_X1 U276 ( .A(n2650), .Z(n2942) );
  BUF_X1 U277 ( .A(n2647), .Z(n2945) );
  BUF_X1 U278 ( .A(n2644), .Z(n2948) );
  BUF_X1 U279 ( .A(n2641), .Z(n2951) );
  BUF_X1 U280 ( .A(n2638), .Z(n2954) );
  BUF_X1 U281 ( .A(n2635), .Z(n2957) );
  BUF_X1 U282 ( .A(n2632), .Z(n2960) );
  BUF_X1 U283 ( .A(n2629), .Z(n2963) );
  BUF_X1 U284 ( .A(n2626), .Z(n2966) );
  BUF_X1 U285 ( .A(n2623), .Z(n2969) );
  BUF_X1 U286 ( .A(n2620), .Z(n2972) );
  BUF_X1 U287 ( .A(n2617), .Z(n2975) );
  BUF_X1 U288 ( .A(n2614), .Z(n2978) );
  BUF_X1 U289 ( .A(n2611), .Z(n2981) );
  BUF_X1 U290 ( .A(n2608), .Z(n2984) );
  BUF_X1 U291 ( .A(n2605), .Z(n2987) );
  BUF_X1 U292 ( .A(n2602), .Z(n2989) );
  BUF_X1 U293 ( .A(n2599), .Z(n2992) );
  BUF_X1 U294 ( .A(n2596), .Z(n2995) );
  BUF_X1 U295 ( .A(n2593), .Z(n2998) );
  BUF_X1 U296 ( .A(n2590), .Z(n3001) );
  BUF_X1 U297 ( .A(n2587), .Z(n3004) );
  BUF_X1 U298 ( .A(n2584), .Z(n3007) );
  BUF_X1 U299 ( .A(n2581), .Z(n3010) );
  BUF_X1 U300 ( .A(n2578), .Z(n3013) );
  BUF_X1 U301 ( .A(n2575), .Z(n3016) );
  BUF_X1 U302 ( .A(n2572), .Z(n3019) );
  BUF_X1 U303 ( .A(n2569), .Z(n3022) );
  BUF_X1 U304 ( .A(n2566), .Z(n3025) );
  BUF_X1 U305 ( .A(n2563), .Z(n3028) );
  BUF_X1 U306 ( .A(n2560), .Z(n3031) );
  BUF_X1 U307 ( .A(n2557), .Z(n3034) );
  BUF_X1 U308 ( .A(n2554), .Z(n3037) );
  BUF_X1 U309 ( .A(n2551), .Z(n3040) );
  BUF_X1 U310 ( .A(n2548), .Z(n3043) );
  BUF_X1 U311 ( .A(n2545), .Z(n3046) );
  BUF_X1 U312 ( .A(n2542), .Z(n3049) );
  BUF_X1 U313 ( .A(n2539), .Z(n3052) );
  BUF_X1 U314 ( .A(n2536), .Z(n3055) );
  BUF_X1 U315 ( .A(n2533), .Z(n3058) );
  BUF_X1 U316 ( .A(n2530), .Z(n3061) );
  BUF_X1 U317 ( .A(n2527), .Z(n3064) );
  BUF_X1 U318 ( .A(n2524), .Z(n3067) );
  BUF_X1 U319 ( .A(n2521), .Z(n3070) );
  BUF_X1 U320 ( .A(n2518), .Z(n3073) );
  BUF_X1 U321 ( .A(n2515), .Z(n3076) );
  BUF_X1 U322 ( .A(n2512), .Z(n3079) );
  BUF_X1 U323 ( .A(n2506), .Z(n3085) );
  BUF_X1 U324 ( .A(n2602), .Z(n2988) );
  BUF_X1 U325 ( .A(n2599), .Z(n2991) );
  BUF_X1 U326 ( .A(n2596), .Z(n2994) );
  BUF_X1 U327 ( .A(n2593), .Z(n2997) );
  BUF_X1 U328 ( .A(n2590), .Z(n3000) );
  BUF_X1 U329 ( .A(n2587), .Z(n3003) );
  BUF_X1 U330 ( .A(n2584), .Z(n3006) );
  BUF_X1 U331 ( .A(n2581), .Z(n3009) );
  BUF_X1 U332 ( .A(n2578), .Z(n3012) );
  BUF_X1 U333 ( .A(n2575), .Z(n3015) );
  BUF_X1 U334 ( .A(n2572), .Z(n3018) );
  BUF_X1 U335 ( .A(n2569), .Z(n3021) );
  BUF_X1 U336 ( .A(n2566), .Z(n3024) );
  BUF_X1 U337 ( .A(n2563), .Z(n3027) );
  BUF_X1 U338 ( .A(n2560), .Z(n3030) );
  BUF_X1 U339 ( .A(n2557), .Z(n3033) );
  BUF_X1 U340 ( .A(n2554), .Z(n3036) );
  BUF_X1 U341 ( .A(n2551), .Z(n3039) );
  BUF_X1 U342 ( .A(n2548), .Z(n3042) );
  BUF_X1 U343 ( .A(n2545), .Z(n3045) );
  BUF_X1 U344 ( .A(n2542), .Z(n3048) );
  BUF_X1 U345 ( .A(n2539), .Z(n3051) );
  BUF_X1 U346 ( .A(n2536), .Z(n3054) );
  BUF_X1 U347 ( .A(n2533), .Z(n3057) );
  BUF_X1 U348 ( .A(n2530), .Z(n3060) );
  BUF_X1 U349 ( .A(n2527), .Z(n3063) );
  BUF_X1 U350 ( .A(n2524), .Z(n3066) );
  BUF_X1 U351 ( .A(n2521), .Z(n3069) );
  BUF_X1 U352 ( .A(n2518), .Z(n3072) );
  BUF_X1 U353 ( .A(n2515), .Z(n3075) );
  BUF_X1 U354 ( .A(n2512), .Z(n3078) );
  BUF_X1 U355 ( .A(n2506), .Z(n3084) );
  BUF_X1 U356 ( .A(n2602), .Z(n2990) );
  BUF_X1 U357 ( .A(n2599), .Z(n2993) );
  BUF_X1 U358 ( .A(n2596), .Z(n2996) );
  BUF_X1 U359 ( .A(n2593), .Z(n2999) );
  BUF_X1 U360 ( .A(n2590), .Z(n3002) );
  BUF_X1 U361 ( .A(n2587), .Z(n3005) );
  BUF_X1 U362 ( .A(n2584), .Z(n3008) );
  BUF_X1 U363 ( .A(n2581), .Z(n3011) );
  BUF_X1 U364 ( .A(n2578), .Z(n3014) );
  BUF_X1 U365 ( .A(n2575), .Z(n3017) );
  BUF_X1 U366 ( .A(n2572), .Z(n3020) );
  BUF_X1 U367 ( .A(n2569), .Z(n3023) );
  BUF_X1 U368 ( .A(n2566), .Z(n3026) );
  BUF_X1 U369 ( .A(n2563), .Z(n3029) );
  BUF_X1 U370 ( .A(n2560), .Z(n3032) );
  BUF_X1 U371 ( .A(n2557), .Z(n3035) );
  BUF_X1 U372 ( .A(n2554), .Z(n3038) );
  BUF_X1 U373 ( .A(n2551), .Z(n3041) );
  BUF_X1 U374 ( .A(n2548), .Z(n3044) );
  BUF_X1 U375 ( .A(n2545), .Z(n3047) );
  BUF_X1 U376 ( .A(n2542), .Z(n3050) );
  BUF_X1 U377 ( .A(n2539), .Z(n3053) );
  BUF_X1 U378 ( .A(n2536), .Z(n3056) );
  BUF_X1 U379 ( .A(n2533), .Z(n3059) );
  BUF_X1 U380 ( .A(n2530), .Z(n3062) );
  BUF_X1 U381 ( .A(n2527), .Z(n3065) );
  BUF_X1 U382 ( .A(n2524), .Z(n3068) );
  BUF_X1 U383 ( .A(n2521), .Z(n3071) );
  BUF_X1 U384 ( .A(n2518), .Z(n3074) );
  BUF_X1 U385 ( .A(n2515), .Z(n3077) );
  BUF_X1 U386 ( .A(n2512), .Z(n3080) );
  BUF_X1 U387 ( .A(n2506), .Z(n3086) );
  AND3_X1 U388 ( .A1(n2303), .A2(n2305), .A3(n3099), .ZN(n2285) );
  AND3_X1 U389 ( .A1(n1677), .A2(n1681), .A3(n3099), .ZN(n1649) );
  OAI21_X1 U390 ( .B1(n526), .B2(n527), .A(n3096), .ZN(n2695) );
  OAI21_X1 U391 ( .B1(n526), .B2(n528), .A(n3095), .ZN(n2692) );
  OAI21_X1 U392 ( .B1(n526), .B2(n529), .A(n3095), .ZN(n2689) );
  OAI21_X1 U393 ( .B1(n526), .B2(n530), .A(n3095), .ZN(n2686) );
  OAI21_X1 U394 ( .B1(n526), .B2(n531), .A(n3095), .ZN(n2683) );
  OAI21_X1 U395 ( .B1(n526), .B2(n532), .A(n3095), .ZN(n2680) );
  OAI21_X1 U396 ( .B1(n526), .B2(n533), .A(n3095), .ZN(n2677) );
  OAI21_X1 U397 ( .B1(n526), .B2(n534), .A(n3095), .ZN(n2674) );
  OAI21_X1 U398 ( .B1(n527), .B2(n536), .A(n3095), .ZN(n2671) );
  OAI21_X1 U399 ( .B1(n528), .B2(n536), .A(n3095), .ZN(n2668) );
  OAI21_X1 U400 ( .B1(n529), .B2(n536), .A(n3095), .ZN(n2665) );
  OAI21_X1 U401 ( .B1(n530), .B2(n536), .A(n3096), .ZN(n2662) );
  OAI21_X1 U402 ( .B1(n531), .B2(n536), .A(n3096), .ZN(n2659) );
  OAI21_X1 U403 ( .B1(n532), .B2(n536), .A(n3096), .ZN(n2656) );
  OAI21_X1 U404 ( .B1(n533), .B2(n536), .A(n3095), .ZN(n2653) );
  OAI21_X1 U405 ( .B1(n534), .B2(n536), .A(n3096), .ZN(n2650) );
  OAI21_X1 U406 ( .B1(n527), .B2(n538), .A(n3096), .ZN(n2647) );
  OAI21_X1 U407 ( .B1(n528), .B2(n538), .A(n3096), .ZN(n2644) );
  OAI21_X1 U408 ( .B1(n529), .B2(n538), .A(n3096), .ZN(n2641) );
  OAI21_X1 U409 ( .B1(n530), .B2(n538), .A(n3096), .ZN(n2638) );
  OAI21_X1 U410 ( .B1(n531), .B2(n538), .A(n3096), .ZN(n2635) );
  OAI21_X1 U411 ( .B1(n532), .B2(n538), .A(n3096), .ZN(n2632) );
  OAI21_X1 U412 ( .B1(n533), .B2(n538), .A(n3097), .ZN(n2629) );
  OAI21_X1 U413 ( .B1(n534), .B2(n538), .A(n3097), .ZN(n2626) );
  OAI21_X1 U414 ( .B1(n527), .B2(n540), .A(n3097), .ZN(n2623) );
  OAI21_X1 U415 ( .B1(n528), .B2(n540), .A(n3097), .ZN(n2620) );
  OAI21_X1 U416 ( .B1(n529), .B2(n540), .A(n3097), .ZN(n2617) );
  OAI21_X1 U417 ( .B1(n530), .B2(n540), .A(n3096), .ZN(n2614) );
  OAI21_X1 U418 ( .B1(n531), .B2(n540), .A(n3097), .ZN(n2611) );
  OAI21_X1 U419 ( .B1(n532), .B2(n540), .A(n3097), .ZN(n2608) );
  OAI21_X1 U420 ( .B1(n533), .B2(n540), .A(n3097), .ZN(n2605) );
  BUF_X1 U421 ( .A(n3094), .Z(n3099) );
  BUF_X1 U422 ( .A(n3093), .Z(n3096) );
  BUF_X1 U423 ( .A(n3093), .Z(n3095) );
  BUF_X1 U424 ( .A(n3093), .Z(n3097) );
  BUF_X1 U425 ( .A(n3094), .Z(n3098) );
  NAND2_X1 U426 ( .A1(n2297), .A2(n2282), .ZN(n1713) );
  NAND2_X1 U427 ( .A1(n2298), .A2(n2282), .ZN(n1712) );
  NAND2_X1 U428 ( .A1(n2297), .A2(n2285), .ZN(n1718) );
  NAND2_X1 U429 ( .A1(n2298), .A2(n2285), .ZN(n1717) );
  NAND2_X1 U430 ( .A1(n2301), .A2(n2282), .ZN(n1723) );
  NAND2_X1 U431 ( .A1(n2302), .A2(n2282), .ZN(n1722) );
  NAND2_X1 U432 ( .A1(n2301), .A2(n2285), .ZN(n1728) );
  NAND2_X1 U433 ( .A1(n2302), .A2(n2285), .ZN(n1727) );
  NAND2_X1 U434 ( .A1(n1668), .A2(n1644), .ZN(n584) );
  NAND2_X1 U435 ( .A1(n1667), .A2(n1644), .ZN(n586) );
  NAND2_X1 U436 ( .A1(n1668), .A2(n1649), .ZN(n591) );
  NAND2_X1 U437 ( .A1(n1667), .A2(n1649), .ZN(n593) );
  NAND2_X1 U438 ( .A1(n1676), .A2(n1644), .ZN(n598) );
  NAND2_X1 U439 ( .A1(n1675), .A2(n1644), .ZN(n600) );
  NAND2_X1 U440 ( .A1(n1676), .A2(n1649), .ZN(n605) );
  NAND2_X1 U441 ( .A1(n1675), .A2(n1649), .ZN(n607) );
  NAND2_X1 U442 ( .A1(n2282), .A2(n2288), .ZN(n1699) );
  NAND2_X1 U443 ( .A1(n2282), .A2(n2289), .ZN(n1698) );
  NAND2_X1 U444 ( .A1(n1644), .A2(n1655), .ZN(n566) );
  NAND2_X1 U445 ( .A1(n1644), .A2(n1654), .ZN(n568) );
  NAND2_X1 U446 ( .A1(n2285), .A2(n2288), .ZN(n1704) );
  NAND2_X1 U447 ( .A1(n2285), .A2(n2289), .ZN(n1703) );
  NAND2_X1 U448 ( .A1(n1649), .A2(n1655), .ZN(n573) );
  NAND2_X1 U449 ( .A1(n1649), .A2(n1654), .ZN(n575) );
  NAND2_X1 U450 ( .A1(n2279), .A2(n2282), .ZN(n1689) );
  NAND2_X1 U451 ( .A1(n2281), .A2(n2282), .ZN(n1688) );
  NAND2_X1 U452 ( .A1(n2279), .A2(n2285), .ZN(n1694) );
  NAND2_X1 U453 ( .A1(n2281), .A2(n2285), .ZN(n1693) );
  NAND2_X1 U454 ( .A1(n1643), .A2(n1644), .ZN(n552) );
  NAND2_X1 U455 ( .A1(n1641), .A2(n1644), .ZN(n554) );
  NAND2_X1 U456 ( .A1(n1643), .A2(n1649), .ZN(n559) );
  NAND2_X1 U457 ( .A1(n1641), .A2(n1649), .ZN(n561) );
  BUF_X1 U458 ( .A(n2503), .Z(n3087) );
  BUF_X1 U459 ( .A(n2503), .Z(n3088) );
  BUF_X1 U460 ( .A(n2500), .Z(n3090) );
  BUF_X1 U461 ( .A(n2500), .Z(n3091) );
  AND2_X1 U462 ( .A1(n2297), .A2(n2280), .ZN(n1716) );
  AND2_X1 U463 ( .A1(n2298), .A2(n2280), .ZN(n1715) );
  AND2_X1 U464 ( .A1(n2297), .A2(n2284), .ZN(n1721) );
  AND2_X1 U465 ( .A1(n2298), .A2(n2284), .ZN(n1720) );
  AND2_X1 U466 ( .A1(n2301), .A2(n2280), .ZN(n1726) );
  AND2_X1 U467 ( .A1(n2302), .A2(n2280), .ZN(n1725) );
  AND2_X1 U468 ( .A1(n2301), .A2(n2284), .ZN(n1731) );
  AND2_X1 U469 ( .A1(n2302), .A2(n2284), .ZN(n1730) );
  AND2_X1 U470 ( .A1(n1668), .A2(n1642), .ZN(n589) );
  AND2_X1 U471 ( .A1(n1667), .A2(n1642), .ZN(n590) );
  AND2_X1 U472 ( .A1(n1668), .A2(n1648), .ZN(n596) );
  AND2_X1 U473 ( .A1(n1667), .A2(n1648), .ZN(n597) );
  AND2_X1 U474 ( .A1(n1676), .A2(n1642), .ZN(n603) );
  AND2_X1 U475 ( .A1(n1675), .A2(n1642), .ZN(n604) );
  AND2_X1 U476 ( .A1(n1676), .A2(n1648), .ZN(n610) );
  AND2_X1 U477 ( .A1(n1675), .A2(n1648), .ZN(n611) );
  BUF_X1 U478 ( .A(n2503), .Z(n3089) );
  BUF_X1 U479 ( .A(n2500), .Z(n3092) );
  AND2_X1 U480 ( .A1(n2284), .A2(n2289), .ZN(n1706) );
  AND2_X1 U481 ( .A1(n1648), .A2(n1655), .ZN(n578) );
  AND2_X1 U482 ( .A1(n1642), .A2(n1655), .ZN(n571) );
  AND2_X1 U483 ( .A1(n1642), .A2(n1654), .ZN(n572) );
  AND2_X1 U484 ( .A1(n2280), .A2(n2288), .ZN(n1702) );
  AND2_X1 U485 ( .A1(n2280), .A2(n2289), .ZN(n1701) );
  AND2_X1 U486 ( .A1(n2279), .A2(n2284), .ZN(n1697) );
  AND2_X1 U487 ( .A1(n2281), .A2(n2284), .ZN(n1696) );
  AND2_X1 U488 ( .A1(n2288), .A2(n2284), .ZN(n1707) );
  AND2_X1 U489 ( .A1(n1643), .A2(n1648), .ZN(n564) );
  AND2_X1 U490 ( .A1(n1641), .A2(n1648), .ZN(n565) );
  AND2_X1 U491 ( .A1(n1654), .A2(n1648), .ZN(n579) );
  AND2_X1 U492 ( .A1(n1643), .A2(n1642), .ZN(n557) );
  AND2_X1 U493 ( .A1(n1641), .A2(n1642), .ZN(n558) );
  AND2_X1 U494 ( .A1(n2279), .A2(n2280), .ZN(n1692) );
  AND2_X1 U495 ( .A1(n2281), .A2(n2280), .ZN(n1691) );
  NAND2_X1 U496 ( .A1(n2272), .A2(n2273), .ZN(N4403) );
  NOR4_X1 U497 ( .A1(n2292), .A2(n2293), .A3(n2294), .A4(n2295), .ZN(n2272) );
  NOR4_X1 U498 ( .A1(n2274), .A2(n2275), .A3(n2276), .A4(n2277), .ZN(n2273) );
  OAI221_X1 U499 ( .B1(n1678), .B2(n2712), .C1(n1679), .C2(n2709), .A(n2304), 
        .ZN(n2292) );
  NAND2_X1 U500 ( .A1(n2254), .A2(n2255), .ZN(N4405) );
  NOR4_X1 U501 ( .A1(n2264), .A2(n2265), .A3(n2266), .A4(n2267), .ZN(n2254) );
  NOR4_X1 U502 ( .A1(n2256), .A2(n2257), .A3(n2258), .A4(n2259), .ZN(n2255) );
  OAI221_X1 U503 ( .B1(n1629), .B2(n2712), .C1(n1630), .C2(n2709), .A(n2271), 
        .ZN(n2264) );
  NAND2_X1 U504 ( .A1(n2236), .A2(n2237), .ZN(N4407) );
  NOR4_X1 U505 ( .A1(n2246), .A2(n2247), .A3(n2248), .A4(n2249), .ZN(n2236) );
  NOR4_X1 U506 ( .A1(n2238), .A2(n2239), .A3(n2240), .A4(n2241), .ZN(n2237) );
  OAI221_X1 U507 ( .B1(n1595), .B2(n2712), .C1(n1596), .C2(n2709), .A(n2253), 
        .ZN(n2246) );
  NAND2_X1 U508 ( .A1(n2218), .A2(n2219), .ZN(N4409) );
  NOR4_X1 U509 ( .A1(n2228), .A2(n2229), .A3(n2230), .A4(n2231), .ZN(n2218) );
  NOR4_X1 U510 ( .A1(n2220), .A2(n2221), .A3(n2222), .A4(n2223), .ZN(n2219) );
  OAI221_X1 U511 ( .B1(n1561), .B2(n2712), .C1(n1562), .C2(n2709), .A(n2235), 
        .ZN(n2228) );
  NAND2_X1 U512 ( .A1(n2200), .A2(n2201), .ZN(N4411) );
  NOR4_X1 U513 ( .A1(n2210), .A2(n2211), .A3(n2212), .A4(n2213), .ZN(n2200) );
  NOR4_X1 U514 ( .A1(n2202), .A2(n2203), .A3(n2204), .A4(n2205), .ZN(n2201) );
  OAI221_X1 U515 ( .B1(n1527), .B2(n2712), .C1(n1528), .C2(n2709), .A(n2217), 
        .ZN(n2210) );
  NAND2_X1 U516 ( .A1(n2182), .A2(n2183), .ZN(N4413) );
  NOR4_X1 U517 ( .A1(n2192), .A2(n2193), .A3(n2194), .A4(n2195), .ZN(n2182) );
  NOR4_X1 U518 ( .A1(n2184), .A2(n2185), .A3(n2186), .A4(n2187), .ZN(n2183) );
  OAI221_X1 U519 ( .B1(n1493), .B2(n2712), .C1(n1494), .C2(n2709), .A(n2199), 
        .ZN(n2192) );
  NAND2_X1 U520 ( .A1(n2164), .A2(n2165), .ZN(N4415) );
  NOR4_X1 U521 ( .A1(n2174), .A2(n2175), .A3(n2176), .A4(n2177), .ZN(n2164) );
  NOR4_X1 U522 ( .A1(n2166), .A2(n2167), .A3(n2168), .A4(n2169), .ZN(n2165) );
  OAI221_X1 U523 ( .B1(n1459), .B2(n2712), .C1(n1460), .C2(n2709), .A(n2181), 
        .ZN(n2174) );
  NAND2_X1 U524 ( .A1(n2146), .A2(n2147), .ZN(N4417) );
  NOR4_X1 U525 ( .A1(n2156), .A2(n2157), .A3(n2158), .A4(n2159), .ZN(n2146) );
  NOR4_X1 U526 ( .A1(n2148), .A2(n2149), .A3(n2150), .A4(n2151), .ZN(n2147) );
  OAI221_X1 U527 ( .B1(n1425), .B2(n2712), .C1(n1426), .C2(n2709), .A(n2163), 
        .ZN(n2156) );
  NAND2_X1 U528 ( .A1(n2128), .A2(n2129), .ZN(N4419) );
  NOR4_X1 U529 ( .A1(n2138), .A2(n2139), .A3(n2140), .A4(n2141), .ZN(n2128) );
  NOR4_X1 U530 ( .A1(n2130), .A2(n2131), .A3(n2132), .A4(n2133), .ZN(n2129) );
  OAI221_X1 U531 ( .B1(n1391), .B2(n2712), .C1(n1392), .C2(n2709), .A(n2145), 
        .ZN(n2138) );
  NAND2_X1 U532 ( .A1(n2110), .A2(n2111), .ZN(N4421) );
  NOR4_X1 U533 ( .A1(n2120), .A2(n2121), .A3(n2122), .A4(n2123), .ZN(n2110) );
  NOR4_X1 U534 ( .A1(n2112), .A2(n2113), .A3(n2114), .A4(n2115), .ZN(n2111) );
  OAI221_X1 U535 ( .B1(n1357), .B2(n2712), .C1(n1358), .C2(n2709), .A(n2127), 
        .ZN(n2120) );
  NAND2_X1 U536 ( .A1(n2092), .A2(n2093), .ZN(N4423) );
  NOR4_X1 U537 ( .A1(n2102), .A2(n2103), .A3(n2104), .A4(n2105), .ZN(n2092) );
  NOR4_X1 U538 ( .A1(n2094), .A2(n2095), .A3(n2096), .A4(n2097), .ZN(n2093) );
  OAI221_X1 U539 ( .B1(n1323), .B2(n2712), .C1(n1324), .C2(n2709), .A(n2109), 
        .ZN(n2102) );
  NAND2_X1 U540 ( .A1(n2074), .A2(n2075), .ZN(N4425) );
  NOR4_X1 U541 ( .A1(n2084), .A2(n2085), .A3(n2086), .A4(n2087), .ZN(n2074) );
  NOR4_X1 U542 ( .A1(n2076), .A2(n2077), .A3(n2078), .A4(n2079), .ZN(n2075) );
  OAI221_X1 U543 ( .B1(n1289), .B2(n2712), .C1(n1290), .C2(n2709), .A(n2091), 
        .ZN(n2084) );
  NAND2_X1 U544 ( .A1(n2056), .A2(n2057), .ZN(N4427) );
  NOR4_X1 U545 ( .A1(n2066), .A2(n2067), .A3(n2068), .A4(n2069), .ZN(n2056) );
  NOR4_X1 U546 ( .A1(n2058), .A2(n2059), .A3(n2060), .A4(n2061), .ZN(n2057) );
  OAI221_X1 U547 ( .B1(n1255), .B2(n2713), .C1(n1256), .C2(n2710), .A(n2073), 
        .ZN(n2066) );
  NAND2_X1 U548 ( .A1(n2038), .A2(n2039), .ZN(N4429) );
  NOR4_X1 U549 ( .A1(n2048), .A2(n2049), .A3(n2050), .A4(n2051), .ZN(n2038) );
  NOR4_X1 U550 ( .A1(n2040), .A2(n2041), .A3(n2042), .A4(n2043), .ZN(n2039) );
  OAI221_X1 U551 ( .B1(n1221), .B2(n2713), .C1(n1222), .C2(n2710), .A(n2055), 
        .ZN(n2048) );
  NAND2_X1 U552 ( .A1(n2020), .A2(n2021), .ZN(N4431) );
  NOR4_X1 U553 ( .A1(n2030), .A2(n2031), .A3(n2032), .A4(n2033), .ZN(n2020) );
  NOR4_X1 U554 ( .A1(n2022), .A2(n2023), .A3(n2024), .A4(n2025), .ZN(n2021) );
  OAI221_X1 U555 ( .B1(n1187), .B2(n2713), .C1(n1188), .C2(n2710), .A(n2037), 
        .ZN(n2030) );
  NAND2_X1 U556 ( .A1(n2002), .A2(n2003), .ZN(N4433) );
  NOR4_X1 U557 ( .A1(n2012), .A2(n2013), .A3(n2014), .A4(n2015), .ZN(n2002) );
  NOR4_X1 U558 ( .A1(n2004), .A2(n2005), .A3(n2006), .A4(n2007), .ZN(n2003) );
  OAI221_X1 U559 ( .B1(n1153), .B2(n2713), .C1(n1154), .C2(n2710), .A(n2019), 
        .ZN(n2012) );
  NAND2_X1 U560 ( .A1(n1984), .A2(n1985), .ZN(N4435) );
  NOR4_X1 U561 ( .A1(n1994), .A2(n1995), .A3(n1996), .A4(n1997), .ZN(n1984) );
  NOR4_X1 U562 ( .A1(n1986), .A2(n1987), .A3(n1988), .A4(n1989), .ZN(n1985) );
  OAI221_X1 U563 ( .B1(n1119), .B2(n2713), .C1(n1120), .C2(n2710), .A(n2001), 
        .ZN(n1994) );
  NAND2_X1 U564 ( .A1(n1966), .A2(n1967), .ZN(N4437) );
  NOR4_X1 U565 ( .A1(n1976), .A2(n1977), .A3(n1978), .A4(n1979), .ZN(n1966) );
  NOR4_X1 U566 ( .A1(n1968), .A2(n1969), .A3(n1970), .A4(n1971), .ZN(n1967) );
  OAI221_X1 U567 ( .B1(n1085), .B2(n2713), .C1(n1086), .C2(n2710), .A(n1983), 
        .ZN(n1976) );
  NAND2_X1 U568 ( .A1(n1948), .A2(n1949), .ZN(N4439) );
  NOR4_X1 U569 ( .A1(n1958), .A2(n1959), .A3(n1960), .A4(n1961), .ZN(n1948) );
  NOR4_X1 U570 ( .A1(n1950), .A2(n1951), .A3(n1952), .A4(n1953), .ZN(n1949) );
  OAI221_X1 U571 ( .B1(n1051), .B2(n2713), .C1(n1052), .C2(n2710), .A(n1965), 
        .ZN(n1958) );
  NAND2_X1 U572 ( .A1(n1930), .A2(n1931), .ZN(N4441) );
  NOR4_X1 U573 ( .A1(n1940), .A2(n1941), .A3(n1942), .A4(n1943), .ZN(n1930) );
  NOR4_X1 U574 ( .A1(n1932), .A2(n1933), .A3(n1934), .A4(n1935), .ZN(n1931) );
  OAI221_X1 U575 ( .B1(n1017), .B2(n2713), .C1(n1018), .C2(n2710), .A(n1947), 
        .ZN(n1940) );
  NAND2_X1 U576 ( .A1(n1912), .A2(n1913), .ZN(N4443) );
  NOR4_X1 U577 ( .A1(n1922), .A2(n1923), .A3(n1924), .A4(n1925), .ZN(n1912) );
  NOR4_X1 U578 ( .A1(n1914), .A2(n1915), .A3(n1916), .A4(n1917), .ZN(n1913) );
  OAI221_X1 U579 ( .B1(n983), .B2(n2713), .C1(n984), .C2(n2710), .A(n1929), 
        .ZN(n1922) );
  NAND2_X1 U580 ( .A1(n1894), .A2(n1895), .ZN(N4445) );
  NOR4_X1 U581 ( .A1(n1904), .A2(n1905), .A3(n1906), .A4(n1907), .ZN(n1894) );
  NOR4_X1 U582 ( .A1(n1896), .A2(n1897), .A3(n1898), .A4(n1899), .ZN(n1895) );
  OAI221_X1 U583 ( .B1(n949), .B2(n2713), .C1(n950), .C2(n2710), .A(n1911), 
        .ZN(n1904) );
  NAND2_X1 U584 ( .A1(n1876), .A2(n1877), .ZN(N4447) );
  NOR4_X1 U585 ( .A1(n1886), .A2(n1887), .A3(n1888), .A4(n1889), .ZN(n1876) );
  NOR4_X1 U586 ( .A1(n1878), .A2(n1879), .A3(n1880), .A4(n1881), .ZN(n1877) );
  OAI221_X1 U587 ( .B1(n915), .B2(n2713), .C1(n916), .C2(n2710), .A(n1893), 
        .ZN(n1886) );
  NAND2_X1 U588 ( .A1(n1858), .A2(n1859), .ZN(N4449) );
  NOR4_X1 U589 ( .A1(n1868), .A2(n1869), .A3(n1870), .A4(n1871), .ZN(n1858) );
  NOR4_X1 U590 ( .A1(n1860), .A2(n1861), .A3(n1862), .A4(n1863), .ZN(n1859) );
  OAI221_X1 U591 ( .B1(n881), .B2(n2713), .C1(n882), .C2(n2710), .A(n1875), 
        .ZN(n1868) );
  NAND2_X1 U592 ( .A1(n1840), .A2(n1841), .ZN(N4451) );
  NOR4_X1 U593 ( .A1(n1850), .A2(n1851), .A3(n1852), .A4(n1853), .ZN(n1840) );
  NOR4_X1 U594 ( .A1(n1842), .A2(n1843), .A3(n1844), .A4(n1845), .ZN(n1841) );
  OAI221_X1 U595 ( .B1(n847), .B2(n2714), .C1(n848), .C2(n2711), .A(n1857), 
        .ZN(n1850) );
  NAND2_X1 U596 ( .A1(n1822), .A2(n1823), .ZN(N4453) );
  NOR4_X1 U597 ( .A1(n1832), .A2(n1833), .A3(n1834), .A4(n1835), .ZN(n1822) );
  NOR4_X1 U598 ( .A1(n1824), .A2(n1825), .A3(n1826), .A4(n1827), .ZN(n1823) );
  OAI221_X1 U599 ( .B1(n813), .B2(n2714), .C1(n814), .C2(n2711), .A(n1839), 
        .ZN(n1832) );
  NAND2_X1 U600 ( .A1(n1804), .A2(n1805), .ZN(N4455) );
  NOR4_X1 U601 ( .A1(n1814), .A2(n1815), .A3(n1816), .A4(n1817), .ZN(n1804) );
  NOR4_X1 U602 ( .A1(n1806), .A2(n1807), .A3(n1808), .A4(n1809), .ZN(n1805) );
  OAI221_X1 U603 ( .B1(n779), .B2(n2714), .C1(n780), .C2(n2711), .A(n1821), 
        .ZN(n1814) );
  NAND2_X1 U604 ( .A1(n1786), .A2(n1787), .ZN(N4457) );
  NOR4_X1 U605 ( .A1(n1796), .A2(n1797), .A3(n1798), .A4(n1799), .ZN(n1786) );
  NOR4_X1 U606 ( .A1(n1788), .A2(n1789), .A3(n1790), .A4(n1791), .ZN(n1787) );
  OAI221_X1 U607 ( .B1(n745), .B2(n2714), .C1(n746), .C2(n2711), .A(n1803), 
        .ZN(n1796) );
  NAND2_X1 U608 ( .A1(n1768), .A2(n1769), .ZN(N4459) );
  NOR4_X1 U609 ( .A1(n1778), .A2(n1779), .A3(n1780), .A4(n1781), .ZN(n1768) );
  NOR4_X1 U610 ( .A1(n1770), .A2(n1771), .A3(n1772), .A4(n1773), .ZN(n1769) );
  OAI221_X1 U611 ( .B1(n711), .B2(n2714), .C1(n712), .C2(n2711), .A(n1785), 
        .ZN(n1778) );
  NAND2_X1 U612 ( .A1(n1750), .A2(n1751), .ZN(N4461) );
  NOR4_X1 U613 ( .A1(n1760), .A2(n1761), .A3(n1762), .A4(n1763), .ZN(n1750) );
  NOR4_X1 U614 ( .A1(n1752), .A2(n1753), .A3(n1754), .A4(n1755), .ZN(n1751) );
  OAI221_X1 U615 ( .B1(n677), .B2(n2714), .C1(n678), .C2(n2711), .A(n1767), 
        .ZN(n1760) );
  NAND2_X1 U616 ( .A1(n1732), .A2(n1733), .ZN(N4463) );
  NOR4_X1 U617 ( .A1(n1742), .A2(n1743), .A3(n1744), .A4(n1745), .ZN(n1732) );
  NOR4_X1 U618 ( .A1(n1734), .A2(n1735), .A3(n1736), .A4(n1737), .ZN(n1733) );
  OAI221_X1 U619 ( .B1(n643), .B2(n2714), .C1(n644), .C2(n2711), .A(n1749), 
        .ZN(n1742) );
  NAND2_X1 U620 ( .A1(n1682), .A2(n1683), .ZN(N4465) );
  NOR4_X1 U621 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(n1682) );
  NOR4_X1 U622 ( .A1(n1684), .A2(n1685), .A3(n1686), .A4(n1687), .ZN(n1683) );
  OAI221_X1 U623 ( .B1(n606), .B2(n2714), .C1(n608), .C2(n2711), .A(n1729), 
        .ZN(n1708) );
  NAND2_X1 U624 ( .A1(n1632), .A2(n1633), .ZN(N4467) );
  NOR4_X1 U625 ( .A1(n1660), .A2(n1661), .A3(n1662), .A4(n1663), .ZN(n1632) );
  NOR4_X1 U626 ( .A1(n1634), .A2(n1635), .A3(n1636), .A4(n1637), .ZN(n1633) );
  OAI221_X1 U627 ( .B1(n2808), .B2(n1678), .C1(n2805), .C2(n1679), .A(n1680), 
        .ZN(n1660) );
  NAND2_X1 U628 ( .A1(n1598), .A2(n1599), .ZN(N4469) );
  NOR4_X1 U629 ( .A1(n1616), .A2(n1617), .A3(n1618), .A4(n1619), .ZN(n1598) );
  NOR4_X1 U630 ( .A1(n1600), .A2(n1601), .A3(n1602), .A4(n1603), .ZN(n1599) );
  OAI221_X1 U631 ( .B1(n2808), .B2(n1629), .C1(n2805), .C2(n1630), .A(n1631), 
        .ZN(n1616) );
  NAND2_X1 U632 ( .A1(n1564), .A2(n1565), .ZN(N4471) );
  NOR4_X1 U633 ( .A1(n1582), .A2(n1583), .A3(n1584), .A4(n1585), .ZN(n1564) );
  NOR4_X1 U634 ( .A1(n1566), .A2(n1567), .A3(n1568), .A4(n1569), .ZN(n1565) );
  OAI221_X1 U635 ( .B1(n2808), .B2(n1595), .C1(n2805), .C2(n1596), .A(n1597), 
        .ZN(n1582) );
  NAND2_X1 U636 ( .A1(n1530), .A2(n1531), .ZN(N4473) );
  NOR4_X1 U637 ( .A1(n1548), .A2(n1549), .A3(n1550), .A4(n1551), .ZN(n1530) );
  NOR4_X1 U638 ( .A1(n1532), .A2(n1533), .A3(n1534), .A4(n1535), .ZN(n1531) );
  OAI221_X1 U639 ( .B1(n2808), .B2(n1561), .C1(n2805), .C2(n1562), .A(n1563), 
        .ZN(n1548) );
  NAND2_X1 U640 ( .A1(n1496), .A2(n1497), .ZN(N4475) );
  NOR4_X1 U641 ( .A1(n1514), .A2(n1515), .A3(n1516), .A4(n1517), .ZN(n1496) );
  NOR4_X1 U642 ( .A1(n1498), .A2(n1499), .A3(n1500), .A4(n1501), .ZN(n1497) );
  OAI221_X1 U643 ( .B1(n2808), .B2(n1527), .C1(n2805), .C2(n1528), .A(n1529), 
        .ZN(n1514) );
  NAND2_X1 U644 ( .A1(n1462), .A2(n1463), .ZN(N4477) );
  NOR4_X1 U645 ( .A1(n1480), .A2(n1481), .A3(n1482), .A4(n1483), .ZN(n1462) );
  NOR4_X1 U646 ( .A1(n1464), .A2(n1465), .A3(n1466), .A4(n1467), .ZN(n1463) );
  OAI221_X1 U647 ( .B1(n2808), .B2(n1493), .C1(n2805), .C2(n1494), .A(n1495), 
        .ZN(n1480) );
  NAND2_X1 U648 ( .A1(n1428), .A2(n1429), .ZN(N4479) );
  NOR4_X1 U649 ( .A1(n1446), .A2(n1447), .A3(n1448), .A4(n1449), .ZN(n1428) );
  NOR4_X1 U650 ( .A1(n1430), .A2(n1431), .A3(n1432), .A4(n1433), .ZN(n1429) );
  OAI221_X1 U651 ( .B1(n2808), .B2(n1459), .C1(n2805), .C2(n1460), .A(n1461), 
        .ZN(n1446) );
  NAND2_X1 U652 ( .A1(n1394), .A2(n1395), .ZN(N4481) );
  NOR4_X1 U653 ( .A1(n1412), .A2(n1413), .A3(n1414), .A4(n1415), .ZN(n1394) );
  NOR4_X1 U654 ( .A1(n1396), .A2(n1397), .A3(n1398), .A4(n1399), .ZN(n1395) );
  OAI221_X1 U655 ( .B1(n2808), .B2(n1425), .C1(n2805), .C2(n1426), .A(n1427), 
        .ZN(n1412) );
  NAND2_X1 U656 ( .A1(n1360), .A2(n1361), .ZN(N4483) );
  NOR4_X1 U657 ( .A1(n1378), .A2(n1379), .A3(n1380), .A4(n1381), .ZN(n1360) );
  NOR4_X1 U658 ( .A1(n1362), .A2(n1363), .A3(n1364), .A4(n1365), .ZN(n1361) );
  OAI221_X1 U659 ( .B1(n2808), .B2(n1391), .C1(n2805), .C2(n1392), .A(n1393), 
        .ZN(n1378) );
  NAND2_X1 U660 ( .A1(n1326), .A2(n1327), .ZN(N4485) );
  NOR4_X1 U661 ( .A1(n1344), .A2(n1345), .A3(n1346), .A4(n1347), .ZN(n1326) );
  NOR4_X1 U662 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1331), .ZN(n1327) );
  OAI221_X1 U663 ( .B1(n2808), .B2(n1357), .C1(n2805), .C2(n1358), .A(n1359), 
        .ZN(n1344) );
  NAND2_X1 U664 ( .A1(n1292), .A2(n1293), .ZN(N4487) );
  NOR4_X1 U665 ( .A1(n1310), .A2(n1311), .A3(n1312), .A4(n1313), .ZN(n1292) );
  NOR4_X1 U666 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1293) );
  OAI221_X1 U667 ( .B1(n2808), .B2(n1323), .C1(n2805), .C2(n1324), .A(n1325), 
        .ZN(n1310) );
  NAND2_X1 U668 ( .A1(n1258), .A2(n1259), .ZN(N4489) );
  NOR4_X1 U669 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1258) );
  NOR4_X1 U670 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1259) );
  OAI221_X1 U671 ( .B1(n2808), .B2(n1289), .C1(n2805), .C2(n1290), .A(n1291), 
        .ZN(n1276) );
  NAND2_X1 U672 ( .A1(n1224), .A2(n1225), .ZN(N4491) );
  NOR4_X1 U673 ( .A1(n1242), .A2(n1243), .A3(n1244), .A4(n1245), .ZN(n1224) );
  NOR4_X1 U674 ( .A1(n1226), .A2(n1227), .A3(n1228), .A4(n1229), .ZN(n1225) );
  OAI221_X1 U675 ( .B1(n2809), .B2(n1255), .C1(n2806), .C2(n1256), .A(n1257), 
        .ZN(n1242) );
  NAND2_X1 U676 ( .A1(n1190), .A2(n1191), .ZN(N4493) );
  NOR4_X1 U677 ( .A1(n1208), .A2(n1209), .A3(n1210), .A4(n1211), .ZN(n1190) );
  NOR4_X1 U678 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n1191) );
  OAI221_X1 U679 ( .B1(n2809), .B2(n1221), .C1(n2806), .C2(n1222), .A(n1223), 
        .ZN(n1208) );
  NAND2_X1 U680 ( .A1(n1156), .A2(n1157), .ZN(N4495) );
  NOR4_X1 U681 ( .A1(n1174), .A2(n1175), .A3(n1176), .A4(n1177), .ZN(n1156) );
  NOR4_X1 U682 ( .A1(n1158), .A2(n1159), .A3(n1160), .A4(n1161), .ZN(n1157) );
  OAI221_X1 U683 ( .B1(n2809), .B2(n1187), .C1(n2806), .C2(n1188), .A(n1189), 
        .ZN(n1174) );
  NAND2_X1 U684 ( .A1(n1122), .A2(n1123), .ZN(N4497) );
  NOR4_X1 U685 ( .A1(n1140), .A2(n1141), .A3(n1142), .A4(n1143), .ZN(n1122) );
  NOR4_X1 U686 ( .A1(n1124), .A2(n1125), .A3(n1126), .A4(n1127), .ZN(n1123) );
  OAI221_X1 U687 ( .B1(n2809), .B2(n1153), .C1(n2806), .C2(n1154), .A(n1155), 
        .ZN(n1140) );
  NAND2_X1 U688 ( .A1(n1088), .A2(n1089), .ZN(N4499) );
  NOR4_X1 U689 ( .A1(n1106), .A2(n1107), .A3(n1108), .A4(n1109), .ZN(n1088) );
  NOR4_X1 U690 ( .A1(n1090), .A2(n1091), .A3(n1092), .A4(n1093), .ZN(n1089) );
  OAI221_X1 U691 ( .B1(n2809), .B2(n1119), .C1(n2806), .C2(n1120), .A(n1121), 
        .ZN(n1106) );
  NAND2_X1 U692 ( .A1(n1054), .A2(n1055), .ZN(N4501) );
  NOR4_X1 U693 ( .A1(n1072), .A2(n1073), .A3(n1074), .A4(n1075), .ZN(n1054) );
  NOR4_X1 U694 ( .A1(n1056), .A2(n1057), .A3(n1058), .A4(n1059), .ZN(n1055) );
  OAI221_X1 U695 ( .B1(n2809), .B2(n1085), .C1(n2806), .C2(n1086), .A(n1087), 
        .ZN(n1072) );
  NAND2_X1 U696 ( .A1(n1020), .A2(n1021), .ZN(N4503) );
  NOR4_X1 U697 ( .A1(n1038), .A2(n1039), .A3(n1040), .A4(n1041), .ZN(n1020) );
  NOR4_X1 U698 ( .A1(n1022), .A2(n1023), .A3(n1024), .A4(n1025), .ZN(n1021) );
  OAI221_X1 U699 ( .B1(n2809), .B2(n1051), .C1(n2806), .C2(n1052), .A(n1053), 
        .ZN(n1038) );
  NAND2_X1 U700 ( .A1(n986), .A2(n987), .ZN(N4505) );
  NOR4_X1 U701 ( .A1(n1004), .A2(n1005), .A3(n1006), .A4(n1007), .ZN(n986) );
  NOR4_X1 U702 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .ZN(n987) );
  OAI221_X1 U703 ( .B1(n2809), .B2(n1017), .C1(n2806), .C2(n1018), .A(n1019), 
        .ZN(n1004) );
  NAND2_X1 U704 ( .A1(n952), .A2(n953), .ZN(N4507) );
  NOR4_X1 U705 ( .A1(n970), .A2(n971), .A3(n972), .A4(n973), .ZN(n952) );
  NOR4_X1 U706 ( .A1(n954), .A2(n955), .A3(n956), .A4(n957), .ZN(n953) );
  OAI221_X1 U707 ( .B1(n2809), .B2(n983), .C1(n2806), .C2(n984), .A(n985), 
        .ZN(n970) );
  NAND2_X1 U708 ( .A1(n918), .A2(n919), .ZN(N4509) );
  NOR4_X1 U709 ( .A1(n936), .A2(n937), .A3(n938), .A4(n939), .ZN(n918) );
  NOR4_X1 U710 ( .A1(n920), .A2(n921), .A3(n922), .A4(n923), .ZN(n919) );
  OAI221_X1 U711 ( .B1(n2809), .B2(n949), .C1(n2806), .C2(n950), .A(n951), 
        .ZN(n936) );
  NAND2_X1 U712 ( .A1(n884), .A2(n885), .ZN(N4511) );
  NOR4_X1 U713 ( .A1(n902), .A2(n903), .A3(n904), .A4(n905), .ZN(n884) );
  NOR4_X1 U714 ( .A1(n886), .A2(n887), .A3(n888), .A4(n889), .ZN(n885) );
  OAI221_X1 U715 ( .B1(n2809), .B2(n915), .C1(n2806), .C2(n916), .A(n917), 
        .ZN(n902) );
  NAND2_X1 U716 ( .A1(n850), .A2(n851), .ZN(N4513) );
  NOR4_X1 U717 ( .A1(n868), .A2(n869), .A3(n870), .A4(n871), .ZN(n850) );
  NOR4_X1 U718 ( .A1(n852), .A2(n853), .A3(n854), .A4(n855), .ZN(n851) );
  OAI221_X1 U719 ( .B1(n2809), .B2(n881), .C1(n2806), .C2(n882), .A(n883), 
        .ZN(n868) );
  NAND2_X1 U720 ( .A1(n816), .A2(n817), .ZN(N4515) );
  NOR4_X1 U721 ( .A1(n834), .A2(n835), .A3(n836), .A4(n837), .ZN(n816) );
  NOR4_X1 U722 ( .A1(n818), .A2(n819), .A3(n820), .A4(n821), .ZN(n817) );
  OAI221_X1 U723 ( .B1(n2810), .B2(n847), .C1(n2807), .C2(n848), .A(n849), 
        .ZN(n834) );
  NAND2_X1 U724 ( .A1(n782), .A2(n783), .ZN(N4517) );
  NOR4_X1 U725 ( .A1(n800), .A2(n801), .A3(n802), .A4(n803), .ZN(n782) );
  NOR4_X1 U726 ( .A1(n784), .A2(n785), .A3(n786), .A4(n787), .ZN(n783) );
  OAI221_X1 U727 ( .B1(n2810), .B2(n813), .C1(n2807), .C2(n814), .A(n815), 
        .ZN(n800) );
  NAND2_X1 U728 ( .A1(n748), .A2(n749), .ZN(N4519) );
  NOR4_X1 U729 ( .A1(n766), .A2(n767), .A3(n768), .A4(n769), .ZN(n748) );
  NOR4_X1 U730 ( .A1(n750), .A2(n751), .A3(n752), .A4(n753), .ZN(n749) );
  OAI221_X1 U731 ( .B1(n2810), .B2(n779), .C1(n2807), .C2(n780), .A(n781), 
        .ZN(n766) );
  NAND2_X1 U732 ( .A1(n714), .A2(n715), .ZN(N4521) );
  NOR4_X1 U733 ( .A1(n732), .A2(n733), .A3(n734), .A4(n735), .ZN(n714) );
  NOR4_X1 U734 ( .A1(n716), .A2(n717), .A3(n718), .A4(n719), .ZN(n715) );
  OAI221_X1 U735 ( .B1(n2810), .B2(n745), .C1(n2807), .C2(n746), .A(n747), 
        .ZN(n732) );
  NAND2_X1 U736 ( .A1(n680), .A2(n681), .ZN(N4523) );
  NOR4_X1 U737 ( .A1(n698), .A2(n699), .A3(n700), .A4(n701), .ZN(n680) );
  NOR4_X1 U738 ( .A1(n682), .A2(n683), .A3(n684), .A4(n685), .ZN(n681) );
  OAI221_X1 U739 ( .B1(n2810), .B2(n711), .C1(n2807), .C2(n712), .A(n713), 
        .ZN(n698) );
  NAND2_X1 U740 ( .A1(n646), .A2(n647), .ZN(N4525) );
  NOR4_X1 U741 ( .A1(n664), .A2(n665), .A3(n666), .A4(n667), .ZN(n646) );
  NOR4_X1 U742 ( .A1(n648), .A2(n649), .A3(n650), .A4(n651), .ZN(n647) );
  OAI221_X1 U743 ( .B1(n2810), .B2(n677), .C1(n2807), .C2(n678), .A(n679), 
        .ZN(n664) );
  NAND2_X1 U744 ( .A1(n612), .A2(n613), .ZN(N4527) );
  NOR4_X1 U745 ( .A1(n630), .A2(n631), .A3(n632), .A4(n633), .ZN(n612) );
  NOR4_X1 U746 ( .A1(n614), .A2(n615), .A3(n616), .A4(n617), .ZN(n613) );
  OAI221_X1 U747 ( .B1(n2810), .B2(n643), .C1(n2807), .C2(n644), .A(n645), 
        .ZN(n630) );
  NAND2_X1 U748 ( .A1(n546), .A2(n547), .ZN(N4529) );
  NOR4_X1 U749 ( .A1(n580), .A2(n581), .A3(n582), .A4(n583), .ZN(n546) );
  NOR4_X1 U750 ( .A1(n548), .A2(n549), .A3(n550), .A4(n551), .ZN(n547) );
  OAI221_X1 U751 ( .B1(n2810), .B2(n606), .C1(n2807), .C2(n608), .A(n609), 
        .ZN(n580) );
  AND2_X1 U752 ( .A1(DATAIN[20]), .A2(n3099), .ZN(n2542) );
  AND2_X1 U753 ( .A1(DATAIN[21]), .A2(n3099), .ZN(n2539) );
  AND2_X1 U754 ( .A1(DATAIN[22]), .A2(n3099), .ZN(n2536) );
  AND2_X1 U755 ( .A1(DATAIN[23]), .A2(n3099), .ZN(n2533) );
  AND2_X1 U756 ( .A1(DATAIN[25]), .A2(n3099), .ZN(n2527) );
  AND2_X1 U757 ( .A1(DATAIN[26]), .A2(n3099), .ZN(n2524) );
  AND2_X1 U758 ( .A1(DATAIN[27]), .A2(n3099), .ZN(n2521) );
  AND2_X1 U759 ( .A1(DATAIN[28]), .A2(n3099), .ZN(n2518) );
  AND2_X1 U760 ( .A1(DATAIN[29]), .A2(n3099), .ZN(n2515) );
  AND2_X1 U761 ( .A1(DATAIN[30]), .A2(n3099), .ZN(n2512) );
  AND2_X1 U762 ( .A1(DATAIN[31]), .A2(n3099), .ZN(n2506) );
  AND2_X1 U763 ( .A1(DATAIN[0]), .A2(n3097), .ZN(n2602) );
  AND2_X1 U764 ( .A1(DATAIN[1]), .A2(n3097), .ZN(n2599) );
  AND2_X1 U765 ( .A1(DATAIN[2]), .A2(n3097), .ZN(n2596) );
  AND2_X1 U766 ( .A1(DATAIN[3]), .A2(n3098), .ZN(n2593) );
  AND2_X1 U767 ( .A1(DATAIN[4]), .A2(n3098), .ZN(n2590) );
  AND2_X1 U768 ( .A1(DATAIN[5]), .A2(n3098), .ZN(n2587) );
  AND2_X1 U769 ( .A1(DATAIN[6]), .A2(n3098), .ZN(n2584) );
  AND2_X1 U770 ( .A1(DATAIN[7]), .A2(n3098), .ZN(n2581) );
  AND2_X1 U771 ( .A1(DATAIN[8]), .A2(n3098), .ZN(n2578) );
  AND2_X1 U772 ( .A1(DATAIN[9]), .A2(n3098), .ZN(n2575) );
  AND2_X1 U773 ( .A1(DATAIN[10]), .A2(n3098), .ZN(n2572) );
  AND2_X1 U774 ( .A1(DATAIN[11]), .A2(n3098), .ZN(n2569) );
  AND2_X1 U775 ( .A1(DATAIN[12]), .A2(n3098), .ZN(n2566) );
  AND2_X1 U776 ( .A1(DATAIN[13]), .A2(n3098), .ZN(n2563) );
  AND2_X1 U777 ( .A1(DATAIN[14]), .A2(n3098), .ZN(n2560) );
  AND2_X1 U778 ( .A1(DATAIN[15]), .A2(n3098), .ZN(n2557) );
  AND2_X1 U779 ( .A1(DATAIN[16]), .A2(n3098), .ZN(n2554) );
  AND2_X1 U780 ( .A1(DATAIN[17]), .A2(n3098), .ZN(n2551) );
  AND2_X1 U781 ( .A1(DATAIN[18]), .A2(n3098), .ZN(n2548) );
  AND2_X1 U782 ( .A1(DATAIN[19]), .A2(n3098), .ZN(n2545) );
  AND2_X1 U783 ( .A1(DATAIN[24]), .A2(n3098), .ZN(n2530) );
  NOR3_X1 U784 ( .A1(n2286), .A2(ADD_RD1[4]), .A3(n2291), .ZN(n2297) );
  NOR3_X1 U785 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n2291), .ZN(n2298) );
  NOR3_X1 U786 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n2286), .ZN(n2301) );
  NOR3_X1 U787 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n2302)
         );
  NOR3_X1 U788 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n1659), .ZN(n1668) );
  NOR3_X1 U789 ( .A1(n1650), .A2(ADD_RD2[4]), .A3(n1659), .ZN(n1667) );
  NOR3_X1 U790 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n1676)
         );
  NOR3_X1 U791 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n1650), .ZN(n1675) );
  AND3_X1 U792 ( .A1(n3099), .A2(n2303), .A3(ADD_RD1[2]), .ZN(n2282) );
  AND3_X1 U793 ( .A1(n3099), .A2(n1677), .A3(ADD_RD2[2]), .ZN(n1644) );
  OAI221_X1 U794 ( .B1(n2894), .B2(n822), .C1(n2891), .C2(n823), .A(n824), 
        .ZN(n821) );
  AOI22_X1 U795 ( .A1(\REGISTERS[30][24] ), .A2(n2888), .B1(
        \REGISTERS[31][24] ), .B2(n2885), .ZN(n824) );
  OAI221_X1 U796 ( .B1(n2846), .B2(n838), .C1(n2843), .C2(n839), .A(n840), 
        .ZN(n837) );
  AOI22_X1 U797 ( .A1(\REGISTERS[14][24] ), .A2(n2840), .B1(
        \REGISTERS[15][24] ), .B2(n2837), .ZN(n840) );
  OAI221_X1 U798 ( .B1(n2894), .B2(n788), .C1(n2891), .C2(n789), .A(n790), 
        .ZN(n787) );
  AOI22_X1 U799 ( .A1(\REGISTERS[30][25] ), .A2(n2888), .B1(
        \REGISTERS[31][25] ), .B2(n2885), .ZN(n790) );
  OAI221_X1 U800 ( .B1(n2846), .B2(n804), .C1(n2843), .C2(n805), .A(n806), 
        .ZN(n803) );
  AOI22_X1 U801 ( .A1(\REGISTERS[14][25] ), .A2(n2840), .B1(
        \REGISTERS[15][25] ), .B2(n2837), .ZN(n806) );
  OAI221_X1 U802 ( .B1(n2894), .B2(n754), .C1(n2891), .C2(n755), .A(n756), 
        .ZN(n753) );
  AOI22_X1 U803 ( .A1(\REGISTERS[30][26] ), .A2(n2888), .B1(
        \REGISTERS[31][26] ), .B2(n2885), .ZN(n756) );
  OAI221_X1 U804 ( .B1(n2846), .B2(n770), .C1(n2843), .C2(n771), .A(n772), 
        .ZN(n769) );
  AOI22_X1 U805 ( .A1(\REGISTERS[14][26] ), .A2(n2840), .B1(
        \REGISTERS[15][26] ), .B2(n2837), .ZN(n772) );
  OAI221_X1 U806 ( .B1(n2894), .B2(n720), .C1(n2891), .C2(n721), .A(n722), 
        .ZN(n719) );
  AOI22_X1 U807 ( .A1(\REGISTERS[30][27] ), .A2(n2888), .B1(
        \REGISTERS[31][27] ), .B2(n2885), .ZN(n722) );
  OAI221_X1 U808 ( .B1(n2846), .B2(n736), .C1(n2843), .C2(n737), .A(n738), 
        .ZN(n735) );
  AOI22_X1 U809 ( .A1(\REGISTERS[14][27] ), .A2(n2840), .B1(
        \REGISTERS[15][27] ), .B2(n2837), .ZN(n738) );
  OAI221_X1 U810 ( .B1(n2894), .B2(n686), .C1(n2891), .C2(n687), .A(n688), 
        .ZN(n685) );
  AOI22_X1 U811 ( .A1(\REGISTERS[30][28] ), .A2(n2888), .B1(
        \REGISTERS[31][28] ), .B2(n2885), .ZN(n688) );
  OAI221_X1 U812 ( .B1(n2846), .B2(n702), .C1(n2843), .C2(n703), .A(n704), 
        .ZN(n701) );
  AOI22_X1 U813 ( .A1(\REGISTERS[14][28] ), .A2(n2840), .B1(
        \REGISTERS[15][28] ), .B2(n2837), .ZN(n704) );
  OAI221_X1 U814 ( .B1(n2894), .B2(n652), .C1(n2891), .C2(n653), .A(n654), 
        .ZN(n651) );
  AOI22_X1 U815 ( .A1(\REGISTERS[30][29] ), .A2(n2888), .B1(
        \REGISTERS[31][29] ), .B2(n2885), .ZN(n654) );
  OAI221_X1 U816 ( .B1(n2846), .B2(n668), .C1(n2843), .C2(n669), .A(n670), 
        .ZN(n667) );
  AOI22_X1 U817 ( .A1(\REGISTERS[14][29] ), .A2(n2840), .B1(
        \REGISTERS[15][29] ), .B2(n2837), .ZN(n670) );
  OAI221_X1 U818 ( .B1(n2894), .B2(n618), .C1(n2891), .C2(n619), .A(n620), 
        .ZN(n617) );
  AOI22_X1 U819 ( .A1(\REGISTERS[30][30] ), .A2(n2888), .B1(
        \REGISTERS[31][30] ), .B2(n2885), .ZN(n620) );
  OAI221_X1 U820 ( .B1(n2846), .B2(n634), .C1(n2843), .C2(n635), .A(n636), 
        .ZN(n633) );
  AOI22_X1 U821 ( .A1(\REGISTERS[14][30] ), .A2(n2840), .B1(
        \REGISTERS[15][30] ), .B2(n2837), .ZN(n636) );
  OAI221_X1 U822 ( .B1(n2894), .B2(n553), .C1(n2891), .C2(n555), .A(n556), 
        .ZN(n551) );
  AOI22_X1 U823 ( .A1(\REGISTERS[30][31] ), .A2(n2888), .B1(
        \REGISTERS[31][31] ), .B2(n2885), .ZN(n556) );
  OAI221_X1 U824 ( .B1(n2846), .B2(n585), .C1(n2843), .C2(n587), .A(n588), 
        .ZN(n583) );
  AOI22_X1 U825 ( .A1(\REGISTERS[14][31] ), .A2(n2840), .B1(
        \REGISTERS[15][31] ), .B2(n2837), .ZN(n588) );
  OAI221_X1 U826 ( .B1(n822), .B2(n2798), .C1(n823), .C2(n2795), .A(n1846), 
        .ZN(n1845) );
  AOI22_X1 U827 ( .A1(n2792), .A2(\REGISTERS[30][24] ), .B1(n2787), .B2(
        \REGISTERS[31][24] ), .ZN(n1846) );
  OAI221_X1 U828 ( .B1(n838), .B2(n2750), .C1(n839), .C2(n2747), .A(n1854), 
        .ZN(n1853) );
  AOI22_X1 U829 ( .A1(n2744), .A2(\REGISTERS[14][24] ), .B1(n2739), .B2(
        \REGISTERS[15][24] ), .ZN(n1854) );
  OAI221_X1 U830 ( .B1(n788), .B2(n2798), .C1(n789), .C2(n2795), .A(n1828), 
        .ZN(n1827) );
  AOI22_X1 U831 ( .A1(n2792), .A2(\REGISTERS[30][25] ), .B1(n2787), .B2(
        \REGISTERS[31][25] ), .ZN(n1828) );
  OAI221_X1 U832 ( .B1(n804), .B2(n2750), .C1(n805), .C2(n2747), .A(n1836), 
        .ZN(n1835) );
  AOI22_X1 U833 ( .A1(n2744), .A2(\REGISTERS[14][25] ), .B1(n2739), .B2(
        \REGISTERS[15][25] ), .ZN(n1836) );
  OAI221_X1 U834 ( .B1(n754), .B2(n2798), .C1(n755), .C2(n2795), .A(n1810), 
        .ZN(n1809) );
  AOI22_X1 U835 ( .A1(n2792), .A2(\REGISTERS[30][26] ), .B1(n2787), .B2(
        \REGISTERS[31][26] ), .ZN(n1810) );
  OAI221_X1 U836 ( .B1(n770), .B2(n2750), .C1(n771), .C2(n2747), .A(n1818), 
        .ZN(n1817) );
  AOI22_X1 U837 ( .A1(n2744), .A2(\REGISTERS[14][26] ), .B1(n2739), .B2(
        \REGISTERS[15][26] ), .ZN(n1818) );
  OAI221_X1 U838 ( .B1(n720), .B2(n2798), .C1(n721), .C2(n2795), .A(n1792), 
        .ZN(n1791) );
  AOI22_X1 U839 ( .A1(n2792), .A2(\REGISTERS[30][27] ), .B1(n2787), .B2(
        \REGISTERS[31][27] ), .ZN(n1792) );
  OAI221_X1 U840 ( .B1(n736), .B2(n2750), .C1(n737), .C2(n2747), .A(n1800), 
        .ZN(n1799) );
  AOI22_X1 U841 ( .A1(n2744), .A2(\REGISTERS[14][27] ), .B1(n2739), .B2(
        \REGISTERS[15][27] ), .ZN(n1800) );
  OAI221_X1 U842 ( .B1(n686), .B2(n2798), .C1(n687), .C2(n2795), .A(n1774), 
        .ZN(n1773) );
  AOI22_X1 U843 ( .A1(n2792), .A2(\REGISTERS[30][28] ), .B1(n2787), .B2(
        \REGISTERS[31][28] ), .ZN(n1774) );
  OAI221_X1 U844 ( .B1(n702), .B2(n2750), .C1(n703), .C2(n2747), .A(n1782), 
        .ZN(n1781) );
  AOI22_X1 U845 ( .A1(n2744), .A2(\REGISTERS[14][28] ), .B1(n2739), .B2(
        \REGISTERS[15][28] ), .ZN(n1782) );
  OAI221_X1 U846 ( .B1(n652), .B2(n2798), .C1(n653), .C2(n2795), .A(n1756), 
        .ZN(n1755) );
  AOI22_X1 U847 ( .A1(n2792), .A2(\REGISTERS[30][29] ), .B1(n2787), .B2(
        \REGISTERS[31][29] ), .ZN(n1756) );
  OAI221_X1 U848 ( .B1(n668), .B2(n2750), .C1(n669), .C2(n2747), .A(n1764), 
        .ZN(n1763) );
  AOI22_X1 U849 ( .A1(n2744), .A2(\REGISTERS[14][29] ), .B1(n2739), .B2(
        \REGISTERS[15][29] ), .ZN(n1764) );
  OAI221_X1 U850 ( .B1(n618), .B2(n2798), .C1(n619), .C2(n2795), .A(n1738), 
        .ZN(n1737) );
  AOI22_X1 U851 ( .A1(n2792), .A2(\REGISTERS[30][30] ), .B1(n2787), .B2(
        \REGISTERS[31][30] ), .ZN(n1738) );
  OAI221_X1 U852 ( .B1(n634), .B2(n2750), .C1(n635), .C2(n2747), .A(n1746), 
        .ZN(n1745) );
  AOI22_X1 U853 ( .A1(n2744), .A2(\REGISTERS[14][30] ), .B1(n2739), .B2(
        \REGISTERS[15][30] ), .ZN(n1746) );
  OAI221_X1 U854 ( .B1(n553), .B2(n2798), .C1(n555), .C2(n2795), .A(n1690), 
        .ZN(n1687) );
  AOI22_X1 U855 ( .A1(n2792), .A2(\REGISTERS[30][31] ), .B1(n2787), .B2(
        \REGISTERS[31][31] ), .ZN(n1690) );
  OAI221_X1 U856 ( .B1(n585), .B2(n2750), .C1(n587), .C2(n2747), .A(n1714), 
        .ZN(n1711) );
  AOI22_X1 U857 ( .A1(n2744), .A2(\REGISTERS[14][31] ), .B1(n2739), .B2(
        \REGISTERS[15][31] ), .ZN(n1714) );
  OAI221_X1 U858 ( .B1(n1638), .B2(n2796), .C1(n1639), .C2(n2793), .A(n2278), 
        .ZN(n2277) );
  AOI22_X1 U859 ( .A1(n2790), .A2(\REGISTERS[30][0] ), .B1(n2789), .B2(
        \REGISTERS[31][0] ), .ZN(n2278) );
  OAI221_X1 U860 ( .B1(n1664), .B2(n2748), .C1(n1665), .C2(n2745), .A(n2296), 
        .ZN(n2295) );
  AOI22_X1 U861 ( .A1(n2742), .A2(\REGISTERS[14][0] ), .B1(n2741), .B2(
        \REGISTERS[15][0] ), .ZN(n2296) );
  OAI221_X1 U862 ( .B1(n1604), .B2(n2796), .C1(n1605), .C2(n2793), .A(n2260), 
        .ZN(n2259) );
  AOI22_X1 U863 ( .A1(n2790), .A2(\REGISTERS[30][1] ), .B1(n2789), .B2(
        \REGISTERS[31][1] ), .ZN(n2260) );
  OAI221_X1 U864 ( .B1(n1620), .B2(n2748), .C1(n1621), .C2(n2745), .A(n2268), 
        .ZN(n2267) );
  AOI22_X1 U865 ( .A1(n2742), .A2(\REGISTERS[14][1] ), .B1(n2741), .B2(
        \REGISTERS[15][1] ), .ZN(n2268) );
  OAI221_X1 U866 ( .B1(n1570), .B2(n2796), .C1(n1571), .C2(n2793), .A(n2242), 
        .ZN(n2241) );
  AOI22_X1 U867 ( .A1(n2790), .A2(\REGISTERS[30][2] ), .B1(n2789), .B2(
        \REGISTERS[31][2] ), .ZN(n2242) );
  OAI221_X1 U868 ( .B1(n1586), .B2(n2748), .C1(n1587), .C2(n2745), .A(n2250), 
        .ZN(n2249) );
  AOI22_X1 U869 ( .A1(n2742), .A2(\REGISTERS[14][2] ), .B1(n2741), .B2(
        \REGISTERS[15][2] ), .ZN(n2250) );
  OAI221_X1 U870 ( .B1(n1536), .B2(n2796), .C1(n1537), .C2(n2793), .A(n2224), 
        .ZN(n2223) );
  AOI22_X1 U871 ( .A1(n2790), .A2(\REGISTERS[30][3] ), .B1(n2789), .B2(
        \REGISTERS[31][3] ), .ZN(n2224) );
  OAI221_X1 U872 ( .B1(n1552), .B2(n2748), .C1(n1553), .C2(n2745), .A(n2232), 
        .ZN(n2231) );
  AOI22_X1 U873 ( .A1(n2742), .A2(\REGISTERS[14][3] ), .B1(n2741), .B2(
        \REGISTERS[15][3] ), .ZN(n2232) );
  OAI221_X1 U874 ( .B1(n1502), .B2(n2796), .C1(n1503), .C2(n2793), .A(n2206), 
        .ZN(n2205) );
  AOI22_X1 U875 ( .A1(n2790), .A2(\REGISTERS[30][4] ), .B1(n2789), .B2(
        \REGISTERS[31][4] ), .ZN(n2206) );
  OAI221_X1 U876 ( .B1(n1518), .B2(n2748), .C1(n1519), .C2(n2745), .A(n2214), 
        .ZN(n2213) );
  AOI22_X1 U877 ( .A1(n2742), .A2(\REGISTERS[14][4] ), .B1(n2741), .B2(
        \REGISTERS[15][4] ), .ZN(n2214) );
  OAI221_X1 U878 ( .B1(n1468), .B2(n2796), .C1(n1469), .C2(n2793), .A(n2188), 
        .ZN(n2187) );
  AOI22_X1 U879 ( .A1(n2790), .A2(\REGISTERS[30][5] ), .B1(n2789), .B2(
        \REGISTERS[31][5] ), .ZN(n2188) );
  OAI221_X1 U880 ( .B1(n1484), .B2(n2748), .C1(n1485), .C2(n2745), .A(n2196), 
        .ZN(n2195) );
  AOI22_X1 U881 ( .A1(n2742), .A2(\REGISTERS[14][5] ), .B1(n2741), .B2(
        \REGISTERS[15][5] ), .ZN(n2196) );
  OAI221_X1 U882 ( .B1(n1434), .B2(n2796), .C1(n1435), .C2(n2793), .A(n2170), 
        .ZN(n2169) );
  AOI22_X1 U883 ( .A1(n2790), .A2(\REGISTERS[30][6] ), .B1(n2789), .B2(
        \REGISTERS[31][6] ), .ZN(n2170) );
  OAI221_X1 U884 ( .B1(n1450), .B2(n2748), .C1(n1451), .C2(n2745), .A(n2178), 
        .ZN(n2177) );
  AOI22_X1 U885 ( .A1(n2742), .A2(\REGISTERS[14][6] ), .B1(n2741), .B2(
        \REGISTERS[15][6] ), .ZN(n2178) );
  OAI221_X1 U886 ( .B1(n1400), .B2(n2796), .C1(n1401), .C2(n2793), .A(n2152), 
        .ZN(n2151) );
  AOI22_X1 U887 ( .A1(n2790), .A2(\REGISTERS[30][7] ), .B1(n2789), .B2(
        \REGISTERS[31][7] ), .ZN(n2152) );
  OAI221_X1 U888 ( .B1(n1416), .B2(n2748), .C1(n1417), .C2(n2745), .A(n2160), 
        .ZN(n2159) );
  AOI22_X1 U889 ( .A1(n2742), .A2(\REGISTERS[14][7] ), .B1(n2741), .B2(
        \REGISTERS[15][7] ), .ZN(n2160) );
  OAI221_X1 U890 ( .B1(n1366), .B2(n2796), .C1(n1367), .C2(n2793), .A(n2134), 
        .ZN(n2133) );
  AOI22_X1 U891 ( .A1(n2790), .A2(\REGISTERS[30][8] ), .B1(n2788), .B2(
        \REGISTERS[31][8] ), .ZN(n2134) );
  OAI221_X1 U892 ( .B1(n1382), .B2(n2748), .C1(n1383), .C2(n2745), .A(n2142), 
        .ZN(n2141) );
  AOI22_X1 U893 ( .A1(n2742), .A2(\REGISTERS[14][8] ), .B1(n2740), .B2(
        \REGISTERS[15][8] ), .ZN(n2142) );
  OAI221_X1 U894 ( .B1(n1332), .B2(n2796), .C1(n1333), .C2(n2793), .A(n2116), 
        .ZN(n2115) );
  AOI22_X1 U895 ( .A1(n2790), .A2(\REGISTERS[30][9] ), .B1(n2788), .B2(
        \REGISTERS[31][9] ), .ZN(n2116) );
  OAI221_X1 U896 ( .B1(n1348), .B2(n2748), .C1(n1349), .C2(n2745), .A(n2124), 
        .ZN(n2123) );
  AOI22_X1 U897 ( .A1(n2742), .A2(\REGISTERS[14][9] ), .B1(n2740), .B2(
        \REGISTERS[15][9] ), .ZN(n2124) );
  OAI221_X1 U898 ( .B1(n1298), .B2(n2796), .C1(n1299), .C2(n2793), .A(n2098), 
        .ZN(n2097) );
  AOI22_X1 U899 ( .A1(n2790), .A2(\REGISTERS[30][10] ), .B1(n2788), .B2(
        \REGISTERS[31][10] ), .ZN(n2098) );
  OAI221_X1 U900 ( .B1(n1314), .B2(n2748), .C1(n1315), .C2(n2745), .A(n2106), 
        .ZN(n2105) );
  AOI22_X1 U901 ( .A1(n2742), .A2(\REGISTERS[14][10] ), .B1(n2740), .B2(
        \REGISTERS[15][10] ), .ZN(n2106) );
  OAI221_X1 U902 ( .B1(n1264), .B2(n2796), .C1(n1265), .C2(n2793), .A(n2080), 
        .ZN(n2079) );
  AOI22_X1 U903 ( .A1(n2790), .A2(\REGISTERS[30][11] ), .B1(n2788), .B2(
        \REGISTERS[31][11] ), .ZN(n2080) );
  OAI221_X1 U904 ( .B1(n1280), .B2(n2748), .C1(n1281), .C2(n2745), .A(n2088), 
        .ZN(n2087) );
  AOI22_X1 U905 ( .A1(n2742), .A2(\REGISTERS[14][11] ), .B1(n2740), .B2(
        \REGISTERS[15][11] ), .ZN(n2088) );
  OAI221_X1 U906 ( .B1(n1230), .B2(n2797), .C1(n1231), .C2(n2794), .A(n2062), 
        .ZN(n2061) );
  AOI22_X1 U907 ( .A1(n2791), .A2(\REGISTERS[30][12] ), .B1(n2788), .B2(
        \REGISTERS[31][12] ), .ZN(n2062) );
  OAI221_X1 U908 ( .B1(n1246), .B2(n2749), .C1(n1247), .C2(n2746), .A(n2070), 
        .ZN(n2069) );
  AOI22_X1 U909 ( .A1(n2743), .A2(\REGISTERS[14][12] ), .B1(n2740), .B2(
        \REGISTERS[15][12] ), .ZN(n2070) );
  OAI221_X1 U910 ( .B1(n1196), .B2(n2797), .C1(n1197), .C2(n2794), .A(n2044), 
        .ZN(n2043) );
  AOI22_X1 U911 ( .A1(n2791), .A2(\REGISTERS[30][13] ), .B1(n2788), .B2(
        \REGISTERS[31][13] ), .ZN(n2044) );
  OAI221_X1 U912 ( .B1(n1212), .B2(n2749), .C1(n1213), .C2(n2746), .A(n2052), 
        .ZN(n2051) );
  AOI22_X1 U913 ( .A1(n2743), .A2(\REGISTERS[14][13] ), .B1(n2740), .B2(
        \REGISTERS[15][13] ), .ZN(n2052) );
  OAI221_X1 U914 ( .B1(n1162), .B2(n2797), .C1(n1163), .C2(n2794), .A(n2026), 
        .ZN(n2025) );
  AOI22_X1 U915 ( .A1(n2791), .A2(\REGISTERS[30][14] ), .B1(n2788), .B2(
        \REGISTERS[31][14] ), .ZN(n2026) );
  OAI221_X1 U916 ( .B1(n1178), .B2(n2749), .C1(n1179), .C2(n2746), .A(n2034), 
        .ZN(n2033) );
  AOI22_X1 U917 ( .A1(n2743), .A2(\REGISTERS[14][14] ), .B1(n2740), .B2(
        \REGISTERS[15][14] ), .ZN(n2034) );
  OAI221_X1 U918 ( .B1(n1128), .B2(n2797), .C1(n1129), .C2(n2794), .A(n2008), 
        .ZN(n2007) );
  AOI22_X1 U919 ( .A1(n2791), .A2(\REGISTERS[30][15] ), .B1(n2788), .B2(
        \REGISTERS[31][15] ), .ZN(n2008) );
  OAI221_X1 U920 ( .B1(n1144), .B2(n2749), .C1(n1145), .C2(n2746), .A(n2016), 
        .ZN(n2015) );
  AOI22_X1 U921 ( .A1(n2743), .A2(\REGISTERS[14][15] ), .B1(n2740), .B2(
        \REGISTERS[15][15] ), .ZN(n2016) );
  OAI221_X1 U922 ( .B1(n1094), .B2(n2797), .C1(n1095), .C2(n2794), .A(n1990), 
        .ZN(n1989) );
  AOI22_X1 U923 ( .A1(n2791), .A2(\REGISTERS[30][16] ), .B1(n2788), .B2(
        \REGISTERS[31][16] ), .ZN(n1990) );
  OAI221_X1 U924 ( .B1(n1110), .B2(n2749), .C1(n1111), .C2(n2746), .A(n1998), 
        .ZN(n1997) );
  AOI22_X1 U925 ( .A1(n2743), .A2(\REGISTERS[14][16] ), .B1(n2740), .B2(
        \REGISTERS[15][16] ), .ZN(n1998) );
  OAI221_X1 U926 ( .B1(n1060), .B2(n2797), .C1(n1061), .C2(n2794), .A(n1972), 
        .ZN(n1971) );
  AOI22_X1 U927 ( .A1(n2791), .A2(\REGISTERS[30][17] ), .B1(n2788), .B2(
        \REGISTERS[31][17] ), .ZN(n1972) );
  OAI221_X1 U928 ( .B1(n1076), .B2(n2749), .C1(n1077), .C2(n2746), .A(n1980), 
        .ZN(n1979) );
  AOI22_X1 U929 ( .A1(n2743), .A2(\REGISTERS[14][17] ), .B1(n2740), .B2(
        \REGISTERS[15][17] ), .ZN(n1980) );
  OAI221_X1 U930 ( .B1(n1026), .B2(n2797), .C1(n1027), .C2(n2794), .A(n1954), 
        .ZN(n1953) );
  AOI22_X1 U931 ( .A1(n2791), .A2(\REGISTERS[30][18] ), .B1(n2788), .B2(
        \REGISTERS[31][18] ), .ZN(n1954) );
  OAI221_X1 U932 ( .B1(n1042), .B2(n2749), .C1(n1043), .C2(n2746), .A(n1962), 
        .ZN(n1961) );
  AOI22_X1 U933 ( .A1(n2743), .A2(\REGISTERS[14][18] ), .B1(n2740), .B2(
        \REGISTERS[15][18] ), .ZN(n1962) );
  OAI221_X1 U934 ( .B1(n992), .B2(n2797), .C1(n993), .C2(n2794), .A(n1936), 
        .ZN(n1935) );
  AOI22_X1 U935 ( .A1(n2791), .A2(\REGISTERS[30][19] ), .B1(n2788), .B2(
        \REGISTERS[31][19] ), .ZN(n1936) );
  OAI221_X1 U936 ( .B1(n1008), .B2(n2749), .C1(n1009), .C2(n2746), .A(n1944), 
        .ZN(n1943) );
  AOI22_X1 U937 ( .A1(n2743), .A2(\REGISTERS[14][19] ), .B1(n2740), .B2(
        \REGISTERS[15][19] ), .ZN(n1944) );
  OAI221_X1 U938 ( .B1(n958), .B2(n2797), .C1(n959), .C2(n2794), .A(n1918), 
        .ZN(n1917) );
  AOI22_X1 U939 ( .A1(n2791), .A2(\REGISTERS[30][20] ), .B1(n2787), .B2(
        \REGISTERS[31][20] ), .ZN(n1918) );
  OAI221_X1 U940 ( .B1(n974), .B2(n2749), .C1(n975), .C2(n2746), .A(n1926), 
        .ZN(n1925) );
  AOI22_X1 U941 ( .A1(n2743), .A2(\REGISTERS[14][20] ), .B1(n2739), .B2(
        \REGISTERS[15][20] ), .ZN(n1926) );
  OAI221_X1 U942 ( .B1(n924), .B2(n2797), .C1(n925), .C2(n2794), .A(n1900), 
        .ZN(n1899) );
  AOI22_X1 U943 ( .A1(n2791), .A2(\REGISTERS[30][21] ), .B1(n2787), .B2(
        \REGISTERS[31][21] ), .ZN(n1900) );
  OAI221_X1 U944 ( .B1(n940), .B2(n2749), .C1(n941), .C2(n2746), .A(n1908), 
        .ZN(n1907) );
  AOI22_X1 U945 ( .A1(n2743), .A2(\REGISTERS[14][21] ), .B1(n2739), .B2(
        \REGISTERS[15][21] ), .ZN(n1908) );
  OAI221_X1 U946 ( .B1(n890), .B2(n2797), .C1(n891), .C2(n2794), .A(n1882), 
        .ZN(n1881) );
  AOI22_X1 U947 ( .A1(n2791), .A2(\REGISTERS[30][22] ), .B1(n2787), .B2(
        \REGISTERS[31][22] ), .ZN(n1882) );
  OAI221_X1 U948 ( .B1(n906), .B2(n2749), .C1(n907), .C2(n2746), .A(n1890), 
        .ZN(n1889) );
  AOI22_X1 U949 ( .A1(n2743), .A2(\REGISTERS[14][22] ), .B1(n2739), .B2(
        \REGISTERS[15][22] ), .ZN(n1890) );
  OAI221_X1 U950 ( .B1(n856), .B2(n2797), .C1(n857), .C2(n2794), .A(n1864), 
        .ZN(n1863) );
  AOI22_X1 U951 ( .A1(n2791), .A2(\REGISTERS[30][23] ), .B1(n2787), .B2(
        \REGISTERS[31][23] ), .ZN(n1864) );
  OAI221_X1 U952 ( .B1(n872), .B2(n2749), .C1(n873), .C2(n2746), .A(n1872), 
        .ZN(n1871) );
  AOI22_X1 U953 ( .A1(n2743), .A2(\REGISTERS[14][23] ), .B1(n2739), .B2(
        \REGISTERS[15][23] ), .ZN(n1872) );
  OAI221_X1 U954 ( .B1(n2892), .B2(n1638), .C1(n2889), .C2(n1639), .A(n1640), 
        .ZN(n1637) );
  AOI22_X1 U955 ( .A1(\REGISTERS[30][0] ), .A2(n2886), .B1(\REGISTERS[31][0] ), 
        .B2(n2883), .ZN(n1640) );
  OAI221_X1 U956 ( .B1(n2844), .B2(n1664), .C1(n2841), .C2(n1665), .A(n1666), 
        .ZN(n1663) );
  AOI22_X1 U957 ( .A1(\REGISTERS[14][0] ), .A2(n2838), .B1(\REGISTERS[15][0] ), 
        .B2(n2835), .ZN(n1666) );
  OAI221_X1 U958 ( .B1(n2892), .B2(n1604), .C1(n2889), .C2(n1605), .A(n1606), 
        .ZN(n1603) );
  AOI22_X1 U959 ( .A1(\REGISTERS[30][1] ), .A2(n2886), .B1(\REGISTERS[31][1] ), 
        .B2(n2883), .ZN(n1606) );
  OAI221_X1 U960 ( .B1(n2844), .B2(n1620), .C1(n2841), .C2(n1621), .A(n1622), 
        .ZN(n1619) );
  AOI22_X1 U961 ( .A1(\REGISTERS[14][1] ), .A2(n2838), .B1(\REGISTERS[15][1] ), 
        .B2(n2835), .ZN(n1622) );
  OAI221_X1 U962 ( .B1(n2892), .B2(n1570), .C1(n2889), .C2(n1571), .A(n1572), 
        .ZN(n1569) );
  AOI22_X1 U963 ( .A1(\REGISTERS[30][2] ), .A2(n2886), .B1(\REGISTERS[31][2] ), 
        .B2(n2883), .ZN(n1572) );
  OAI221_X1 U964 ( .B1(n2844), .B2(n1586), .C1(n2841), .C2(n1587), .A(n1588), 
        .ZN(n1585) );
  AOI22_X1 U965 ( .A1(\REGISTERS[14][2] ), .A2(n2838), .B1(\REGISTERS[15][2] ), 
        .B2(n2835), .ZN(n1588) );
  OAI221_X1 U966 ( .B1(n2892), .B2(n1536), .C1(n2889), .C2(n1537), .A(n1538), 
        .ZN(n1535) );
  AOI22_X1 U967 ( .A1(\REGISTERS[30][3] ), .A2(n2886), .B1(\REGISTERS[31][3] ), 
        .B2(n2883), .ZN(n1538) );
  OAI221_X1 U968 ( .B1(n2844), .B2(n1552), .C1(n2841), .C2(n1553), .A(n1554), 
        .ZN(n1551) );
  AOI22_X1 U969 ( .A1(\REGISTERS[14][3] ), .A2(n2838), .B1(\REGISTERS[15][3] ), 
        .B2(n2835), .ZN(n1554) );
  OAI221_X1 U970 ( .B1(n2892), .B2(n1502), .C1(n2889), .C2(n1503), .A(n1504), 
        .ZN(n1501) );
  AOI22_X1 U971 ( .A1(\REGISTERS[30][4] ), .A2(n2886), .B1(\REGISTERS[31][4] ), 
        .B2(n2883), .ZN(n1504) );
  OAI221_X1 U972 ( .B1(n2844), .B2(n1518), .C1(n2841), .C2(n1519), .A(n1520), 
        .ZN(n1517) );
  AOI22_X1 U973 ( .A1(\REGISTERS[14][4] ), .A2(n2838), .B1(\REGISTERS[15][4] ), 
        .B2(n2835), .ZN(n1520) );
  OAI221_X1 U974 ( .B1(n2892), .B2(n1468), .C1(n2889), .C2(n1469), .A(n1470), 
        .ZN(n1467) );
  AOI22_X1 U975 ( .A1(\REGISTERS[30][5] ), .A2(n2886), .B1(\REGISTERS[31][5] ), 
        .B2(n2883), .ZN(n1470) );
  OAI221_X1 U976 ( .B1(n2844), .B2(n1484), .C1(n2841), .C2(n1485), .A(n1486), 
        .ZN(n1483) );
  AOI22_X1 U977 ( .A1(\REGISTERS[14][5] ), .A2(n2838), .B1(\REGISTERS[15][5] ), 
        .B2(n2835), .ZN(n1486) );
  OAI221_X1 U978 ( .B1(n2892), .B2(n1434), .C1(n2889), .C2(n1435), .A(n1436), 
        .ZN(n1433) );
  AOI22_X1 U979 ( .A1(\REGISTERS[30][6] ), .A2(n2886), .B1(\REGISTERS[31][6] ), 
        .B2(n2883), .ZN(n1436) );
  OAI221_X1 U980 ( .B1(n2844), .B2(n1450), .C1(n2841), .C2(n1451), .A(n1452), 
        .ZN(n1449) );
  AOI22_X1 U981 ( .A1(\REGISTERS[14][6] ), .A2(n2838), .B1(\REGISTERS[15][6] ), 
        .B2(n2835), .ZN(n1452) );
  OAI221_X1 U982 ( .B1(n2892), .B2(n1400), .C1(n2889), .C2(n1401), .A(n1402), 
        .ZN(n1399) );
  AOI22_X1 U983 ( .A1(\REGISTERS[30][7] ), .A2(n2886), .B1(\REGISTERS[31][7] ), 
        .B2(n2883), .ZN(n1402) );
  OAI221_X1 U984 ( .B1(n2844), .B2(n1416), .C1(n2841), .C2(n1417), .A(n1418), 
        .ZN(n1415) );
  AOI22_X1 U985 ( .A1(\REGISTERS[14][7] ), .A2(n2838), .B1(\REGISTERS[15][7] ), 
        .B2(n2835), .ZN(n1418) );
  OAI221_X1 U986 ( .B1(n2892), .B2(n1366), .C1(n2889), .C2(n1367), .A(n1368), 
        .ZN(n1365) );
  AOI22_X1 U987 ( .A1(\REGISTERS[30][8] ), .A2(n2886), .B1(\REGISTERS[31][8] ), 
        .B2(n2883), .ZN(n1368) );
  OAI221_X1 U988 ( .B1(n2844), .B2(n1382), .C1(n2841), .C2(n1383), .A(n1384), 
        .ZN(n1381) );
  AOI22_X1 U989 ( .A1(\REGISTERS[14][8] ), .A2(n2838), .B1(\REGISTERS[15][8] ), 
        .B2(n2835), .ZN(n1384) );
  OAI221_X1 U990 ( .B1(n2892), .B2(n1332), .C1(n2889), .C2(n1333), .A(n1334), 
        .ZN(n1331) );
  AOI22_X1 U991 ( .A1(\REGISTERS[30][9] ), .A2(n2886), .B1(\REGISTERS[31][9] ), 
        .B2(n2883), .ZN(n1334) );
  OAI221_X1 U992 ( .B1(n2844), .B2(n1348), .C1(n2841), .C2(n1349), .A(n1350), 
        .ZN(n1347) );
  AOI22_X1 U993 ( .A1(\REGISTERS[14][9] ), .A2(n2838), .B1(\REGISTERS[15][9] ), 
        .B2(n2835), .ZN(n1350) );
  OAI221_X1 U994 ( .B1(n2892), .B2(n1298), .C1(n2889), .C2(n1299), .A(n1300), 
        .ZN(n1297) );
  AOI22_X1 U995 ( .A1(\REGISTERS[30][10] ), .A2(n2886), .B1(
        \REGISTERS[31][10] ), .B2(n2883), .ZN(n1300) );
  OAI221_X1 U996 ( .B1(n2844), .B2(n1314), .C1(n2841), .C2(n1315), .A(n1316), 
        .ZN(n1313) );
  AOI22_X1 U997 ( .A1(\REGISTERS[14][10] ), .A2(n2838), .B1(
        \REGISTERS[15][10] ), .B2(n2835), .ZN(n1316) );
  OAI221_X1 U998 ( .B1(n2892), .B2(n1264), .C1(n2889), .C2(n1265), .A(n1266), 
        .ZN(n1263) );
  AOI22_X1 U999 ( .A1(\REGISTERS[30][11] ), .A2(n2886), .B1(
        \REGISTERS[31][11] ), .B2(n2883), .ZN(n1266) );
  OAI221_X1 U1000 ( .B1(n2844), .B2(n1280), .C1(n2841), .C2(n1281), .A(n1282), 
        .ZN(n1279) );
  AOI22_X1 U1001 ( .A1(\REGISTERS[14][11] ), .A2(n2838), .B1(
        \REGISTERS[15][11] ), .B2(n2835), .ZN(n1282) );
  OAI221_X1 U1002 ( .B1(n2893), .B2(n1230), .C1(n2890), .C2(n1231), .A(n1232), 
        .ZN(n1229) );
  AOI22_X1 U1003 ( .A1(\REGISTERS[30][12] ), .A2(n2887), .B1(
        \REGISTERS[31][12] ), .B2(n2884), .ZN(n1232) );
  OAI221_X1 U1004 ( .B1(n2845), .B2(n1246), .C1(n2842), .C2(n1247), .A(n1248), 
        .ZN(n1245) );
  AOI22_X1 U1005 ( .A1(\REGISTERS[14][12] ), .A2(n2839), .B1(
        \REGISTERS[15][12] ), .B2(n2836), .ZN(n1248) );
  OAI221_X1 U1006 ( .B1(n2893), .B2(n1196), .C1(n2890), .C2(n1197), .A(n1198), 
        .ZN(n1195) );
  AOI22_X1 U1007 ( .A1(\REGISTERS[30][13] ), .A2(n2887), .B1(
        \REGISTERS[31][13] ), .B2(n2884), .ZN(n1198) );
  OAI221_X1 U1008 ( .B1(n2845), .B2(n1212), .C1(n2842), .C2(n1213), .A(n1214), 
        .ZN(n1211) );
  AOI22_X1 U1009 ( .A1(\REGISTERS[14][13] ), .A2(n2839), .B1(
        \REGISTERS[15][13] ), .B2(n2836), .ZN(n1214) );
  OAI221_X1 U1010 ( .B1(n2893), .B2(n1162), .C1(n2890), .C2(n1163), .A(n1164), 
        .ZN(n1161) );
  AOI22_X1 U1011 ( .A1(\REGISTERS[30][14] ), .A2(n2887), .B1(
        \REGISTERS[31][14] ), .B2(n2884), .ZN(n1164) );
  OAI221_X1 U1012 ( .B1(n2845), .B2(n1178), .C1(n2842), .C2(n1179), .A(n1180), 
        .ZN(n1177) );
  AOI22_X1 U1013 ( .A1(\REGISTERS[14][14] ), .A2(n2839), .B1(
        \REGISTERS[15][14] ), .B2(n2836), .ZN(n1180) );
  OAI221_X1 U1014 ( .B1(n2893), .B2(n1128), .C1(n2890), .C2(n1129), .A(n1130), 
        .ZN(n1127) );
  AOI22_X1 U1015 ( .A1(\REGISTERS[30][15] ), .A2(n2887), .B1(
        \REGISTERS[31][15] ), .B2(n2884), .ZN(n1130) );
  OAI221_X1 U1016 ( .B1(n2845), .B2(n1144), .C1(n2842), .C2(n1145), .A(n1146), 
        .ZN(n1143) );
  AOI22_X1 U1017 ( .A1(\REGISTERS[14][15] ), .A2(n2839), .B1(
        \REGISTERS[15][15] ), .B2(n2836), .ZN(n1146) );
  OAI221_X1 U1018 ( .B1(n2893), .B2(n1094), .C1(n2890), .C2(n1095), .A(n1096), 
        .ZN(n1093) );
  AOI22_X1 U1019 ( .A1(\REGISTERS[30][16] ), .A2(n2887), .B1(
        \REGISTERS[31][16] ), .B2(n2884), .ZN(n1096) );
  OAI221_X1 U1020 ( .B1(n2845), .B2(n1110), .C1(n2842), .C2(n1111), .A(n1112), 
        .ZN(n1109) );
  AOI22_X1 U1021 ( .A1(\REGISTERS[14][16] ), .A2(n2839), .B1(
        \REGISTERS[15][16] ), .B2(n2836), .ZN(n1112) );
  OAI221_X1 U1022 ( .B1(n2893), .B2(n1060), .C1(n2890), .C2(n1061), .A(n1062), 
        .ZN(n1059) );
  AOI22_X1 U1023 ( .A1(\REGISTERS[30][17] ), .A2(n2887), .B1(
        \REGISTERS[31][17] ), .B2(n2884), .ZN(n1062) );
  OAI221_X1 U1024 ( .B1(n2845), .B2(n1076), .C1(n2842), .C2(n1077), .A(n1078), 
        .ZN(n1075) );
  AOI22_X1 U1025 ( .A1(\REGISTERS[14][17] ), .A2(n2839), .B1(
        \REGISTERS[15][17] ), .B2(n2836), .ZN(n1078) );
  OAI221_X1 U1026 ( .B1(n2893), .B2(n1026), .C1(n2890), .C2(n1027), .A(n1028), 
        .ZN(n1025) );
  AOI22_X1 U1027 ( .A1(\REGISTERS[30][18] ), .A2(n2887), .B1(
        \REGISTERS[31][18] ), .B2(n2884), .ZN(n1028) );
  OAI221_X1 U1028 ( .B1(n2845), .B2(n1042), .C1(n2842), .C2(n1043), .A(n1044), 
        .ZN(n1041) );
  AOI22_X1 U1029 ( .A1(\REGISTERS[14][18] ), .A2(n2839), .B1(
        \REGISTERS[15][18] ), .B2(n2836), .ZN(n1044) );
  OAI221_X1 U1030 ( .B1(n2893), .B2(n992), .C1(n2890), .C2(n993), .A(n994), 
        .ZN(n991) );
  AOI22_X1 U1031 ( .A1(\REGISTERS[30][19] ), .A2(n2887), .B1(
        \REGISTERS[31][19] ), .B2(n2884), .ZN(n994) );
  OAI221_X1 U1032 ( .B1(n2845), .B2(n1008), .C1(n2842), .C2(n1009), .A(n1010), 
        .ZN(n1007) );
  AOI22_X1 U1033 ( .A1(\REGISTERS[14][19] ), .A2(n2839), .B1(
        \REGISTERS[15][19] ), .B2(n2836), .ZN(n1010) );
  OAI221_X1 U1034 ( .B1(n2893), .B2(n958), .C1(n2890), .C2(n959), .A(n960), 
        .ZN(n957) );
  AOI22_X1 U1035 ( .A1(\REGISTERS[30][20] ), .A2(n2887), .B1(
        \REGISTERS[31][20] ), .B2(n2884), .ZN(n960) );
  OAI221_X1 U1036 ( .B1(n2845), .B2(n974), .C1(n2842), .C2(n975), .A(n976), 
        .ZN(n973) );
  AOI22_X1 U1037 ( .A1(\REGISTERS[14][20] ), .A2(n2839), .B1(
        \REGISTERS[15][20] ), .B2(n2836), .ZN(n976) );
  OAI221_X1 U1038 ( .B1(n2893), .B2(n924), .C1(n2890), .C2(n925), .A(n926), 
        .ZN(n923) );
  AOI22_X1 U1039 ( .A1(\REGISTERS[30][21] ), .A2(n2887), .B1(
        \REGISTERS[31][21] ), .B2(n2884), .ZN(n926) );
  OAI221_X1 U1040 ( .B1(n2845), .B2(n940), .C1(n2842), .C2(n941), .A(n942), 
        .ZN(n939) );
  AOI22_X1 U1041 ( .A1(\REGISTERS[14][21] ), .A2(n2839), .B1(
        \REGISTERS[15][21] ), .B2(n2836), .ZN(n942) );
  OAI221_X1 U1042 ( .B1(n2893), .B2(n890), .C1(n2890), .C2(n891), .A(n892), 
        .ZN(n889) );
  AOI22_X1 U1043 ( .A1(\REGISTERS[30][22] ), .A2(n2887), .B1(
        \REGISTERS[31][22] ), .B2(n2884), .ZN(n892) );
  OAI221_X1 U1044 ( .B1(n2845), .B2(n906), .C1(n2842), .C2(n907), .A(n908), 
        .ZN(n905) );
  AOI22_X1 U1045 ( .A1(\REGISTERS[14][22] ), .A2(n2839), .B1(
        \REGISTERS[15][22] ), .B2(n2836), .ZN(n908) );
  OAI221_X1 U1046 ( .B1(n2893), .B2(n856), .C1(n2890), .C2(n857), .A(n858), 
        .ZN(n855) );
  AOI22_X1 U1047 ( .A1(\REGISTERS[30][23] ), .A2(n2887), .B1(
        \REGISTERS[31][23] ), .B2(n2884), .ZN(n858) );
  OAI221_X1 U1048 ( .B1(n2845), .B2(n872), .C1(n2842), .C2(n873), .A(n874), 
        .ZN(n871) );
  AOI22_X1 U1049 ( .A1(\REGISTERS[14][23] ), .A2(n2839), .B1(
        \REGISTERS[15][23] ), .B2(n2836), .ZN(n874) );
  OAI221_X1 U1050 ( .B1(n2882), .B2(n825), .C1(n2879), .C2(n826), .A(n827), 
        .ZN(n820) );
  AOI22_X1 U1051 ( .A1(\REGISTERS[26][24] ), .A2(n2876), .B1(
        \REGISTERS[27][24] ), .B2(n2873), .ZN(n827) );
  OAI221_X1 U1052 ( .B1(n2834), .B2(n841), .C1(n2831), .C2(n842), .A(n843), 
        .ZN(n836) );
  AOI22_X1 U1053 ( .A1(\REGISTERS[10][24] ), .A2(n2828), .B1(
        \REGISTERS[11][24] ), .B2(n2825), .ZN(n843) );
  OAI221_X1 U1054 ( .B1(n2882), .B2(n791), .C1(n2879), .C2(n792), .A(n793), 
        .ZN(n786) );
  AOI22_X1 U1055 ( .A1(\REGISTERS[26][25] ), .A2(n2876), .B1(
        \REGISTERS[27][25] ), .B2(n2873), .ZN(n793) );
  OAI221_X1 U1056 ( .B1(n2834), .B2(n807), .C1(n2831), .C2(n808), .A(n809), 
        .ZN(n802) );
  AOI22_X1 U1057 ( .A1(\REGISTERS[10][25] ), .A2(n2828), .B1(
        \REGISTERS[11][25] ), .B2(n2825), .ZN(n809) );
  OAI221_X1 U1058 ( .B1(n2882), .B2(n757), .C1(n2879), .C2(n758), .A(n759), 
        .ZN(n752) );
  AOI22_X1 U1059 ( .A1(\REGISTERS[26][26] ), .A2(n2876), .B1(
        \REGISTERS[27][26] ), .B2(n2873), .ZN(n759) );
  OAI221_X1 U1060 ( .B1(n2834), .B2(n773), .C1(n2831), .C2(n774), .A(n775), 
        .ZN(n768) );
  AOI22_X1 U1061 ( .A1(\REGISTERS[10][26] ), .A2(n2828), .B1(
        \REGISTERS[11][26] ), .B2(n2825), .ZN(n775) );
  OAI221_X1 U1062 ( .B1(n2882), .B2(n723), .C1(n2879), .C2(n724), .A(n725), 
        .ZN(n718) );
  AOI22_X1 U1063 ( .A1(\REGISTERS[26][27] ), .A2(n2876), .B1(
        \REGISTERS[27][27] ), .B2(n2873), .ZN(n725) );
  OAI221_X1 U1064 ( .B1(n2834), .B2(n739), .C1(n2831), .C2(n740), .A(n741), 
        .ZN(n734) );
  AOI22_X1 U1065 ( .A1(\REGISTERS[10][27] ), .A2(n2828), .B1(
        \REGISTERS[11][27] ), .B2(n2825), .ZN(n741) );
  OAI221_X1 U1066 ( .B1(n2882), .B2(n689), .C1(n2879), .C2(n690), .A(n691), 
        .ZN(n684) );
  AOI22_X1 U1067 ( .A1(\REGISTERS[26][28] ), .A2(n2876), .B1(
        \REGISTERS[27][28] ), .B2(n2873), .ZN(n691) );
  OAI221_X1 U1068 ( .B1(n2834), .B2(n705), .C1(n2831), .C2(n706), .A(n707), 
        .ZN(n700) );
  AOI22_X1 U1069 ( .A1(\REGISTERS[10][28] ), .A2(n2828), .B1(
        \REGISTERS[11][28] ), .B2(n2825), .ZN(n707) );
  OAI221_X1 U1070 ( .B1(n2882), .B2(n655), .C1(n2879), .C2(n656), .A(n657), 
        .ZN(n650) );
  AOI22_X1 U1071 ( .A1(\REGISTERS[26][29] ), .A2(n2876), .B1(
        \REGISTERS[27][29] ), .B2(n2873), .ZN(n657) );
  OAI221_X1 U1072 ( .B1(n2834), .B2(n671), .C1(n2831), .C2(n672), .A(n673), 
        .ZN(n666) );
  AOI22_X1 U1073 ( .A1(\REGISTERS[10][29] ), .A2(n2828), .B1(
        \REGISTERS[11][29] ), .B2(n2825), .ZN(n673) );
  OAI221_X1 U1074 ( .B1(n2882), .B2(n621), .C1(n2879), .C2(n622), .A(n623), 
        .ZN(n616) );
  AOI22_X1 U1075 ( .A1(\REGISTERS[26][30] ), .A2(n2876), .B1(
        \REGISTERS[27][30] ), .B2(n2873), .ZN(n623) );
  OAI221_X1 U1076 ( .B1(n2834), .B2(n637), .C1(n2831), .C2(n638), .A(n639), 
        .ZN(n632) );
  AOI22_X1 U1077 ( .A1(\REGISTERS[10][30] ), .A2(n2828), .B1(
        \REGISTERS[11][30] ), .B2(n2825), .ZN(n639) );
  OAI221_X1 U1078 ( .B1(n2882), .B2(n560), .C1(n2879), .C2(n562), .A(n563), 
        .ZN(n550) );
  AOI22_X1 U1079 ( .A1(\REGISTERS[26][31] ), .A2(n2876), .B1(
        \REGISTERS[27][31] ), .B2(n2873), .ZN(n563) );
  OAI221_X1 U1080 ( .B1(n2834), .B2(n592), .C1(n2831), .C2(n594), .A(n595), 
        .ZN(n582) );
  AOI22_X1 U1081 ( .A1(\REGISTERS[10][31] ), .A2(n2828), .B1(
        \REGISTERS[11][31] ), .B2(n2825), .ZN(n595) );
  OAI221_X1 U1082 ( .B1(n825), .B2(n2786), .C1(n826), .C2(n2783), .A(n1847), 
        .ZN(n1844) );
  AOI22_X1 U1083 ( .A1(n2780), .A2(\REGISTERS[26][24] ), .B1(n2775), .B2(
        \REGISTERS[27][24] ), .ZN(n1847) );
  OAI221_X1 U1084 ( .B1(n841), .B2(n2738), .C1(n842), .C2(n2735), .A(n1855), 
        .ZN(n1852) );
  AOI22_X1 U1085 ( .A1(n2732), .A2(\REGISTERS[10][24] ), .B1(n2727), .B2(
        \REGISTERS[11][24] ), .ZN(n1855) );
  OAI221_X1 U1086 ( .B1(n791), .B2(n2786), .C1(n792), .C2(n2783), .A(n1829), 
        .ZN(n1826) );
  AOI22_X1 U1087 ( .A1(n2780), .A2(\REGISTERS[26][25] ), .B1(n2775), .B2(
        \REGISTERS[27][25] ), .ZN(n1829) );
  OAI221_X1 U1088 ( .B1(n807), .B2(n2738), .C1(n808), .C2(n2735), .A(n1837), 
        .ZN(n1834) );
  AOI22_X1 U1089 ( .A1(n2732), .A2(\REGISTERS[10][25] ), .B1(n2727), .B2(
        \REGISTERS[11][25] ), .ZN(n1837) );
  OAI221_X1 U1090 ( .B1(n757), .B2(n2786), .C1(n758), .C2(n2783), .A(n1811), 
        .ZN(n1808) );
  AOI22_X1 U1091 ( .A1(n2780), .A2(\REGISTERS[26][26] ), .B1(n2775), .B2(
        \REGISTERS[27][26] ), .ZN(n1811) );
  OAI221_X1 U1092 ( .B1(n773), .B2(n2738), .C1(n774), .C2(n2735), .A(n1819), 
        .ZN(n1816) );
  AOI22_X1 U1093 ( .A1(n2732), .A2(\REGISTERS[10][26] ), .B1(n2727), .B2(
        \REGISTERS[11][26] ), .ZN(n1819) );
  OAI221_X1 U1094 ( .B1(n723), .B2(n2786), .C1(n724), .C2(n2783), .A(n1793), 
        .ZN(n1790) );
  AOI22_X1 U1095 ( .A1(n2780), .A2(\REGISTERS[26][27] ), .B1(n2775), .B2(
        \REGISTERS[27][27] ), .ZN(n1793) );
  OAI221_X1 U1096 ( .B1(n739), .B2(n2738), .C1(n740), .C2(n2735), .A(n1801), 
        .ZN(n1798) );
  AOI22_X1 U1097 ( .A1(n2732), .A2(\REGISTERS[10][27] ), .B1(n2727), .B2(
        \REGISTERS[11][27] ), .ZN(n1801) );
  OAI221_X1 U1098 ( .B1(n689), .B2(n2786), .C1(n690), .C2(n2783), .A(n1775), 
        .ZN(n1772) );
  AOI22_X1 U1099 ( .A1(n2780), .A2(\REGISTERS[26][28] ), .B1(n2775), .B2(
        \REGISTERS[27][28] ), .ZN(n1775) );
  OAI221_X1 U1100 ( .B1(n705), .B2(n2738), .C1(n706), .C2(n2735), .A(n1783), 
        .ZN(n1780) );
  AOI22_X1 U1101 ( .A1(n2732), .A2(\REGISTERS[10][28] ), .B1(n2727), .B2(
        \REGISTERS[11][28] ), .ZN(n1783) );
  OAI221_X1 U1102 ( .B1(n655), .B2(n2786), .C1(n656), .C2(n2783), .A(n1757), 
        .ZN(n1754) );
  AOI22_X1 U1103 ( .A1(n2780), .A2(\REGISTERS[26][29] ), .B1(n2775), .B2(
        \REGISTERS[27][29] ), .ZN(n1757) );
  OAI221_X1 U1104 ( .B1(n671), .B2(n2738), .C1(n672), .C2(n2735), .A(n1765), 
        .ZN(n1762) );
  AOI22_X1 U1105 ( .A1(n2732), .A2(\REGISTERS[10][29] ), .B1(n2727), .B2(
        \REGISTERS[11][29] ), .ZN(n1765) );
  OAI221_X1 U1106 ( .B1(n621), .B2(n2786), .C1(n622), .C2(n2783), .A(n1739), 
        .ZN(n1736) );
  AOI22_X1 U1107 ( .A1(n2780), .A2(\REGISTERS[26][30] ), .B1(n2775), .B2(
        \REGISTERS[27][30] ), .ZN(n1739) );
  OAI221_X1 U1108 ( .B1(n637), .B2(n2738), .C1(n638), .C2(n2735), .A(n1747), 
        .ZN(n1744) );
  AOI22_X1 U1109 ( .A1(n2732), .A2(\REGISTERS[10][30] ), .B1(n2727), .B2(
        \REGISTERS[11][30] ), .ZN(n1747) );
  OAI221_X1 U1110 ( .B1(n560), .B2(n2786), .C1(n562), .C2(n2783), .A(n1695), 
        .ZN(n1686) );
  AOI22_X1 U1111 ( .A1(n2780), .A2(\REGISTERS[26][31] ), .B1(n2775), .B2(
        \REGISTERS[27][31] ), .ZN(n1695) );
  OAI221_X1 U1112 ( .B1(n592), .B2(n2738), .C1(n594), .C2(n2735), .A(n1719), 
        .ZN(n1710) );
  AOI22_X1 U1113 ( .A1(n2732), .A2(\REGISTERS[10][31] ), .B1(n2727), .B2(
        \REGISTERS[11][31] ), .ZN(n1719) );
  OAI221_X1 U1114 ( .B1(n1645), .B2(n2784), .C1(n1646), .C2(n2781), .A(n2283), 
        .ZN(n2276) );
  AOI22_X1 U1115 ( .A1(n2778), .A2(\REGISTERS[26][0] ), .B1(n2777), .B2(
        \REGISTERS[27][0] ), .ZN(n2283) );
  OAI221_X1 U1116 ( .B1(n1669), .B2(n2736), .C1(n1670), .C2(n2733), .A(n2299), 
        .ZN(n2294) );
  AOI22_X1 U1117 ( .A1(n2730), .A2(\REGISTERS[10][0] ), .B1(n2729), .B2(
        \REGISTERS[11][0] ), .ZN(n2299) );
  OAI221_X1 U1118 ( .B1(n1607), .B2(n2784), .C1(n1608), .C2(n2781), .A(n2261), 
        .ZN(n2258) );
  AOI22_X1 U1119 ( .A1(n2778), .A2(\REGISTERS[26][1] ), .B1(n2777), .B2(
        \REGISTERS[27][1] ), .ZN(n2261) );
  OAI221_X1 U1120 ( .B1(n1623), .B2(n2736), .C1(n1624), .C2(n2733), .A(n2269), 
        .ZN(n2266) );
  AOI22_X1 U1121 ( .A1(n2730), .A2(\REGISTERS[10][1] ), .B1(n2729), .B2(
        \REGISTERS[11][1] ), .ZN(n2269) );
  OAI221_X1 U1122 ( .B1(n1573), .B2(n2784), .C1(n1574), .C2(n2781), .A(n2243), 
        .ZN(n2240) );
  AOI22_X1 U1123 ( .A1(n2778), .A2(\REGISTERS[26][2] ), .B1(n2777), .B2(
        \REGISTERS[27][2] ), .ZN(n2243) );
  OAI221_X1 U1124 ( .B1(n1589), .B2(n2736), .C1(n1590), .C2(n2733), .A(n2251), 
        .ZN(n2248) );
  AOI22_X1 U1125 ( .A1(n2730), .A2(\REGISTERS[10][2] ), .B1(n2729), .B2(
        \REGISTERS[11][2] ), .ZN(n2251) );
  OAI221_X1 U1126 ( .B1(n1539), .B2(n2784), .C1(n1540), .C2(n2781), .A(n2225), 
        .ZN(n2222) );
  AOI22_X1 U1127 ( .A1(n2778), .A2(\REGISTERS[26][3] ), .B1(n2777), .B2(
        \REGISTERS[27][3] ), .ZN(n2225) );
  OAI221_X1 U1128 ( .B1(n1555), .B2(n2736), .C1(n1556), .C2(n2733), .A(n2233), 
        .ZN(n2230) );
  AOI22_X1 U1129 ( .A1(n2730), .A2(\REGISTERS[10][3] ), .B1(n2729), .B2(
        \REGISTERS[11][3] ), .ZN(n2233) );
  OAI221_X1 U1130 ( .B1(n1505), .B2(n2784), .C1(n1506), .C2(n2781), .A(n2207), 
        .ZN(n2204) );
  AOI22_X1 U1131 ( .A1(n2778), .A2(\REGISTERS[26][4] ), .B1(n2777), .B2(
        \REGISTERS[27][4] ), .ZN(n2207) );
  OAI221_X1 U1132 ( .B1(n1521), .B2(n2736), .C1(n1522), .C2(n2733), .A(n2215), 
        .ZN(n2212) );
  AOI22_X1 U1133 ( .A1(n2730), .A2(\REGISTERS[10][4] ), .B1(n2729), .B2(
        \REGISTERS[11][4] ), .ZN(n2215) );
  OAI221_X1 U1134 ( .B1(n1471), .B2(n2784), .C1(n1472), .C2(n2781), .A(n2189), 
        .ZN(n2186) );
  AOI22_X1 U1135 ( .A1(n2778), .A2(\REGISTERS[26][5] ), .B1(n2777), .B2(
        \REGISTERS[27][5] ), .ZN(n2189) );
  OAI221_X1 U1136 ( .B1(n1487), .B2(n2736), .C1(n1488), .C2(n2733), .A(n2197), 
        .ZN(n2194) );
  AOI22_X1 U1137 ( .A1(n2730), .A2(\REGISTERS[10][5] ), .B1(n2729), .B2(
        \REGISTERS[11][5] ), .ZN(n2197) );
  OAI221_X1 U1138 ( .B1(n1437), .B2(n2784), .C1(n1438), .C2(n2781), .A(n2171), 
        .ZN(n2168) );
  AOI22_X1 U1139 ( .A1(n2778), .A2(\REGISTERS[26][6] ), .B1(n2777), .B2(
        \REGISTERS[27][6] ), .ZN(n2171) );
  OAI221_X1 U1140 ( .B1(n1453), .B2(n2736), .C1(n1454), .C2(n2733), .A(n2179), 
        .ZN(n2176) );
  AOI22_X1 U1141 ( .A1(n2730), .A2(\REGISTERS[10][6] ), .B1(n2729), .B2(
        \REGISTERS[11][6] ), .ZN(n2179) );
  OAI221_X1 U1142 ( .B1(n1403), .B2(n2784), .C1(n1404), .C2(n2781), .A(n2153), 
        .ZN(n2150) );
  AOI22_X1 U1143 ( .A1(n2778), .A2(\REGISTERS[26][7] ), .B1(n2777), .B2(
        \REGISTERS[27][7] ), .ZN(n2153) );
  OAI221_X1 U1144 ( .B1(n1419), .B2(n2736), .C1(n1420), .C2(n2733), .A(n2161), 
        .ZN(n2158) );
  AOI22_X1 U1145 ( .A1(n2730), .A2(\REGISTERS[10][7] ), .B1(n2729), .B2(
        \REGISTERS[11][7] ), .ZN(n2161) );
  OAI221_X1 U1146 ( .B1(n1369), .B2(n2784), .C1(n1370), .C2(n2781), .A(n2135), 
        .ZN(n2132) );
  AOI22_X1 U1147 ( .A1(n2778), .A2(\REGISTERS[26][8] ), .B1(n2776), .B2(
        \REGISTERS[27][8] ), .ZN(n2135) );
  OAI221_X1 U1148 ( .B1(n1385), .B2(n2736), .C1(n1386), .C2(n2733), .A(n2143), 
        .ZN(n2140) );
  AOI22_X1 U1149 ( .A1(n2730), .A2(\REGISTERS[10][8] ), .B1(n2728), .B2(
        \REGISTERS[11][8] ), .ZN(n2143) );
  OAI221_X1 U1150 ( .B1(n1335), .B2(n2784), .C1(n1336), .C2(n2781), .A(n2117), 
        .ZN(n2114) );
  AOI22_X1 U1151 ( .A1(n2778), .A2(\REGISTERS[26][9] ), .B1(n2776), .B2(
        \REGISTERS[27][9] ), .ZN(n2117) );
  OAI221_X1 U1152 ( .B1(n1351), .B2(n2736), .C1(n1352), .C2(n2733), .A(n2125), 
        .ZN(n2122) );
  AOI22_X1 U1153 ( .A1(n2730), .A2(\REGISTERS[10][9] ), .B1(n2728), .B2(
        \REGISTERS[11][9] ), .ZN(n2125) );
  OAI221_X1 U1154 ( .B1(n1301), .B2(n2784), .C1(n1302), .C2(n2781), .A(n2099), 
        .ZN(n2096) );
  AOI22_X1 U1155 ( .A1(n2778), .A2(\REGISTERS[26][10] ), .B1(n2776), .B2(
        \REGISTERS[27][10] ), .ZN(n2099) );
  OAI221_X1 U1156 ( .B1(n1317), .B2(n2736), .C1(n1318), .C2(n2733), .A(n2107), 
        .ZN(n2104) );
  AOI22_X1 U1157 ( .A1(n2730), .A2(\REGISTERS[10][10] ), .B1(n2728), .B2(
        \REGISTERS[11][10] ), .ZN(n2107) );
  OAI221_X1 U1158 ( .B1(n1267), .B2(n2784), .C1(n1268), .C2(n2781), .A(n2081), 
        .ZN(n2078) );
  AOI22_X1 U1159 ( .A1(n2778), .A2(\REGISTERS[26][11] ), .B1(n2776), .B2(
        \REGISTERS[27][11] ), .ZN(n2081) );
  OAI221_X1 U1160 ( .B1(n1283), .B2(n2736), .C1(n1284), .C2(n2733), .A(n2089), 
        .ZN(n2086) );
  AOI22_X1 U1161 ( .A1(n2730), .A2(\REGISTERS[10][11] ), .B1(n2728), .B2(
        \REGISTERS[11][11] ), .ZN(n2089) );
  OAI221_X1 U1162 ( .B1(n1233), .B2(n2785), .C1(n1234), .C2(n2782), .A(n2063), 
        .ZN(n2060) );
  AOI22_X1 U1163 ( .A1(n2779), .A2(\REGISTERS[26][12] ), .B1(n2776), .B2(
        \REGISTERS[27][12] ), .ZN(n2063) );
  OAI221_X1 U1164 ( .B1(n1249), .B2(n2737), .C1(n1250), .C2(n2734), .A(n2071), 
        .ZN(n2068) );
  AOI22_X1 U1165 ( .A1(n2731), .A2(\REGISTERS[10][12] ), .B1(n2728), .B2(
        \REGISTERS[11][12] ), .ZN(n2071) );
  OAI221_X1 U1166 ( .B1(n1199), .B2(n2785), .C1(n1200), .C2(n2782), .A(n2045), 
        .ZN(n2042) );
  AOI22_X1 U1167 ( .A1(n2779), .A2(\REGISTERS[26][13] ), .B1(n2776), .B2(
        \REGISTERS[27][13] ), .ZN(n2045) );
  OAI221_X1 U1168 ( .B1(n1215), .B2(n2737), .C1(n1216), .C2(n2734), .A(n2053), 
        .ZN(n2050) );
  AOI22_X1 U1169 ( .A1(n2731), .A2(\REGISTERS[10][13] ), .B1(n2728), .B2(
        \REGISTERS[11][13] ), .ZN(n2053) );
  OAI221_X1 U1170 ( .B1(n1165), .B2(n2785), .C1(n1166), .C2(n2782), .A(n2027), 
        .ZN(n2024) );
  AOI22_X1 U1171 ( .A1(n2779), .A2(\REGISTERS[26][14] ), .B1(n2776), .B2(
        \REGISTERS[27][14] ), .ZN(n2027) );
  OAI221_X1 U1172 ( .B1(n1181), .B2(n2737), .C1(n1182), .C2(n2734), .A(n2035), 
        .ZN(n2032) );
  AOI22_X1 U1173 ( .A1(n2731), .A2(\REGISTERS[10][14] ), .B1(n2728), .B2(
        \REGISTERS[11][14] ), .ZN(n2035) );
  OAI221_X1 U1174 ( .B1(n1131), .B2(n2785), .C1(n1132), .C2(n2782), .A(n2009), 
        .ZN(n2006) );
  AOI22_X1 U1175 ( .A1(n2779), .A2(\REGISTERS[26][15] ), .B1(n2776), .B2(
        \REGISTERS[27][15] ), .ZN(n2009) );
  OAI221_X1 U1176 ( .B1(n1147), .B2(n2737), .C1(n1148), .C2(n2734), .A(n2017), 
        .ZN(n2014) );
  AOI22_X1 U1177 ( .A1(n2731), .A2(\REGISTERS[10][15] ), .B1(n2728), .B2(
        \REGISTERS[11][15] ), .ZN(n2017) );
  OAI221_X1 U1178 ( .B1(n1097), .B2(n2785), .C1(n1098), .C2(n2782), .A(n1991), 
        .ZN(n1988) );
  AOI22_X1 U1179 ( .A1(n2779), .A2(\REGISTERS[26][16] ), .B1(n2776), .B2(
        \REGISTERS[27][16] ), .ZN(n1991) );
  OAI221_X1 U1180 ( .B1(n1113), .B2(n2737), .C1(n1114), .C2(n2734), .A(n1999), 
        .ZN(n1996) );
  AOI22_X1 U1181 ( .A1(n2731), .A2(\REGISTERS[10][16] ), .B1(n2728), .B2(
        \REGISTERS[11][16] ), .ZN(n1999) );
  OAI221_X1 U1182 ( .B1(n1063), .B2(n2785), .C1(n1064), .C2(n2782), .A(n1973), 
        .ZN(n1970) );
  AOI22_X1 U1183 ( .A1(n2779), .A2(\REGISTERS[26][17] ), .B1(n2776), .B2(
        \REGISTERS[27][17] ), .ZN(n1973) );
  OAI221_X1 U1184 ( .B1(n1079), .B2(n2737), .C1(n1080), .C2(n2734), .A(n1981), 
        .ZN(n1978) );
  AOI22_X1 U1185 ( .A1(n2731), .A2(\REGISTERS[10][17] ), .B1(n2728), .B2(
        \REGISTERS[11][17] ), .ZN(n1981) );
  OAI221_X1 U1186 ( .B1(n1029), .B2(n2785), .C1(n1030), .C2(n2782), .A(n1955), 
        .ZN(n1952) );
  AOI22_X1 U1187 ( .A1(n2779), .A2(\REGISTERS[26][18] ), .B1(n2776), .B2(
        \REGISTERS[27][18] ), .ZN(n1955) );
  OAI221_X1 U1188 ( .B1(n1045), .B2(n2737), .C1(n1046), .C2(n2734), .A(n1963), 
        .ZN(n1960) );
  AOI22_X1 U1189 ( .A1(n2731), .A2(\REGISTERS[10][18] ), .B1(n2728), .B2(
        \REGISTERS[11][18] ), .ZN(n1963) );
  OAI221_X1 U1190 ( .B1(n995), .B2(n2785), .C1(n996), .C2(n2782), .A(n1937), 
        .ZN(n1934) );
  AOI22_X1 U1191 ( .A1(n2779), .A2(\REGISTERS[26][19] ), .B1(n2776), .B2(
        \REGISTERS[27][19] ), .ZN(n1937) );
  OAI221_X1 U1192 ( .B1(n1011), .B2(n2737), .C1(n1012), .C2(n2734), .A(n1945), 
        .ZN(n1942) );
  AOI22_X1 U1193 ( .A1(n2731), .A2(\REGISTERS[10][19] ), .B1(n2728), .B2(
        \REGISTERS[11][19] ), .ZN(n1945) );
  OAI221_X1 U1194 ( .B1(n961), .B2(n2785), .C1(n962), .C2(n2782), .A(n1919), 
        .ZN(n1916) );
  AOI22_X1 U1195 ( .A1(n2779), .A2(\REGISTERS[26][20] ), .B1(n2775), .B2(
        \REGISTERS[27][20] ), .ZN(n1919) );
  OAI221_X1 U1196 ( .B1(n977), .B2(n2737), .C1(n978), .C2(n2734), .A(n1927), 
        .ZN(n1924) );
  AOI22_X1 U1197 ( .A1(n2731), .A2(\REGISTERS[10][20] ), .B1(n2727), .B2(
        \REGISTERS[11][20] ), .ZN(n1927) );
  OAI221_X1 U1198 ( .B1(n927), .B2(n2785), .C1(n928), .C2(n2782), .A(n1901), 
        .ZN(n1898) );
  AOI22_X1 U1199 ( .A1(n2779), .A2(\REGISTERS[26][21] ), .B1(n2775), .B2(
        \REGISTERS[27][21] ), .ZN(n1901) );
  OAI221_X1 U1200 ( .B1(n943), .B2(n2737), .C1(n944), .C2(n2734), .A(n1909), 
        .ZN(n1906) );
  AOI22_X1 U1201 ( .A1(n2731), .A2(\REGISTERS[10][21] ), .B1(n2727), .B2(
        \REGISTERS[11][21] ), .ZN(n1909) );
  OAI221_X1 U1202 ( .B1(n893), .B2(n2785), .C1(n894), .C2(n2782), .A(n1883), 
        .ZN(n1880) );
  AOI22_X1 U1203 ( .A1(n2779), .A2(\REGISTERS[26][22] ), .B1(n2775), .B2(
        \REGISTERS[27][22] ), .ZN(n1883) );
  OAI221_X1 U1204 ( .B1(n909), .B2(n2737), .C1(n910), .C2(n2734), .A(n1891), 
        .ZN(n1888) );
  AOI22_X1 U1205 ( .A1(n2731), .A2(\REGISTERS[10][22] ), .B1(n2727), .B2(
        \REGISTERS[11][22] ), .ZN(n1891) );
  OAI221_X1 U1206 ( .B1(n859), .B2(n2785), .C1(n860), .C2(n2782), .A(n1865), 
        .ZN(n1862) );
  AOI22_X1 U1207 ( .A1(n2779), .A2(\REGISTERS[26][23] ), .B1(n2775), .B2(
        \REGISTERS[27][23] ), .ZN(n1865) );
  OAI221_X1 U1208 ( .B1(n875), .B2(n2737), .C1(n876), .C2(n2734), .A(n1873), 
        .ZN(n1870) );
  AOI22_X1 U1209 ( .A1(n2731), .A2(\REGISTERS[10][23] ), .B1(n2727), .B2(
        \REGISTERS[11][23] ), .ZN(n1873) );
  OAI221_X1 U1210 ( .B1(n2880), .B2(n1645), .C1(n2877), .C2(n1646), .A(n1647), 
        .ZN(n1636) );
  AOI22_X1 U1211 ( .A1(\REGISTERS[26][0] ), .A2(n2874), .B1(\REGISTERS[27][0] ), .B2(n2871), .ZN(n1647) );
  OAI221_X1 U1212 ( .B1(n2832), .B2(n1669), .C1(n2829), .C2(n1670), .A(n1671), 
        .ZN(n1662) );
  AOI22_X1 U1213 ( .A1(\REGISTERS[10][0] ), .A2(n2826), .B1(\REGISTERS[11][0] ), .B2(n2823), .ZN(n1671) );
  OAI221_X1 U1214 ( .B1(n2880), .B2(n1607), .C1(n2877), .C2(n1608), .A(n1609), 
        .ZN(n1602) );
  AOI22_X1 U1215 ( .A1(\REGISTERS[26][1] ), .A2(n2874), .B1(\REGISTERS[27][1] ), .B2(n2871), .ZN(n1609) );
  OAI221_X1 U1216 ( .B1(n2832), .B2(n1623), .C1(n2829), .C2(n1624), .A(n1625), 
        .ZN(n1618) );
  AOI22_X1 U1217 ( .A1(\REGISTERS[10][1] ), .A2(n2826), .B1(\REGISTERS[11][1] ), .B2(n2823), .ZN(n1625) );
  OAI221_X1 U1218 ( .B1(n2880), .B2(n1573), .C1(n2877), .C2(n1574), .A(n1575), 
        .ZN(n1568) );
  AOI22_X1 U1219 ( .A1(\REGISTERS[26][2] ), .A2(n2874), .B1(\REGISTERS[27][2] ), .B2(n2871), .ZN(n1575) );
  OAI221_X1 U1220 ( .B1(n2832), .B2(n1589), .C1(n2829), .C2(n1590), .A(n1591), 
        .ZN(n1584) );
  AOI22_X1 U1221 ( .A1(\REGISTERS[10][2] ), .A2(n2826), .B1(\REGISTERS[11][2] ), .B2(n2823), .ZN(n1591) );
  OAI221_X1 U1222 ( .B1(n2880), .B2(n1539), .C1(n2877), .C2(n1540), .A(n1541), 
        .ZN(n1534) );
  AOI22_X1 U1223 ( .A1(\REGISTERS[26][3] ), .A2(n2874), .B1(\REGISTERS[27][3] ), .B2(n2871), .ZN(n1541) );
  OAI221_X1 U1224 ( .B1(n2832), .B2(n1555), .C1(n2829), .C2(n1556), .A(n1557), 
        .ZN(n1550) );
  AOI22_X1 U1225 ( .A1(\REGISTERS[10][3] ), .A2(n2826), .B1(\REGISTERS[11][3] ), .B2(n2823), .ZN(n1557) );
  OAI221_X1 U1226 ( .B1(n2880), .B2(n1505), .C1(n2877), .C2(n1506), .A(n1507), 
        .ZN(n1500) );
  AOI22_X1 U1227 ( .A1(\REGISTERS[26][4] ), .A2(n2874), .B1(\REGISTERS[27][4] ), .B2(n2871), .ZN(n1507) );
  OAI221_X1 U1228 ( .B1(n2832), .B2(n1521), .C1(n2829), .C2(n1522), .A(n1523), 
        .ZN(n1516) );
  AOI22_X1 U1229 ( .A1(\REGISTERS[10][4] ), .A2(n2826), .B1(\REGISTERS[11][4] ), .B2(n2823), .ZN(n1523) );
  OAI221_X1 U1230 ( .B1(n2880), .B2(n1471), .C1(n2877), .C2(n1472), .A(n1473), 
        .ZN(n1466) );
  AOI22_X1 U1231 ( .A1(\REGISTERS[26][5] ), .A2(n2874), .B1(\REGISTERS[27][5] ), .B2(n2871), .ZN(n1473) );
  OAI221_X1 U1232 ( .B1(n2832), .B2(n1487), .C1(n2829), .C2(n1488), .A(n1489), 
        .ZN(n1482) );
  AOI22_X1 U1233 ( .A1(\REGISTERS[10][5] ), .A2(n2826), .B1(\REGISTERS[11][5] ), .B2(n2823), .ZN(n1489) );
  OAI221_X1 U1234 ( .B1(n2880), .B2(n1437), .C1(n2877), .C2(n1438), .A(n1439), 
        .ZN(n1432) );
  AOI22_X1 U1235 ( .A1(\REGISTERS[26][6] ), .A2(n2874), .B1(\REGISTERS[27][6] ), .B2(n2871), .ZN(n1439) );
  OAI221_X1 U1236 ( .B1(n2832), .B2(n1453), .C1(n2829), .C2(n1454), .A(n1455), 
        .ZN(n1448) );
  AOI22_X1 U1237 ( .A1(\REGISTERS[10][6] ), .A2(n2826), .B1(\REGISTERS[11][6] ), .B2(n2823), .ZN(n1455) );
  OAI221_X1 U1238 ( .B1(n2880), .B2(n1403), .C1(n2877), .C2(n1404), .A(n1405), 
        .ZN(n1398) );
  AOI22_X1 U1239 ( .A1(\REGISTERS[26][7] ), .A2(n2874), .B1(\REGISTERS[27][7] ), .B2(n2871), .ZN(n1405) );
  OAI221_X1 U1240 ( .B1(n2832), .B2(n1419), .C1(n2829), .C2(n1420), .A(n1421), 
        .ZN(n1414) );
  AOI22_X1 U1241 ( .A1(\REGISTERS[10][7] ), .A2(n2826), .B1(\REGISTERS[11][7] ), .B2(n2823), .ZN(n1421) );
  OAI221_X1 U1242 ( .B1(n2880), .B2(n1369), .C1(n2877), .C2(n1370), .A(n1371), 
        .ZN(n1364) );
  AOI22_X1 U1243 ( .A1(\REGISTERS[26][8] ), .A2(n2874), .B1(\REGISTERS[27][8] ), .B2(n2871), .ZN(n1371) );
  OAI221_X1 U1244 ( .B1(n2832), .B2(n1385), .C1(n2829), .C2(n1386), .A(n1387), 
        .ZN(n1380) );
  AOI22_X1 U1245 ( .A1(\REGISTERS[10][8] ), .A2(n2826), .B1(\REGISTERS[11][8] ), .B2(n2823), .ZN(n1387) );
  OAI221_X1 U1246 ( .B1(n2880), .B2(n1335), .C1(n2877), .C2(n1336), .A(n1337), 
        .ZN(n1330) );
  AOI22_X1 U1247 ( .A1(\REGISTERS[26][9] ), .A2(n2874), .B1(\REGISTERS[27][9] ), .B2(n2871), .ZN(n1337) );
  OAI221_X1 U1248 ( .B1(n2832), .B2(n1351), .C1(n2829), .C2(n1352), .A(n1353), 
        .ZN(n1346) );
  AOI22_X1 U1249 ( .A1(\REGISTERS[10][9] ), .A2(n2826), .B1(\REGISTERS[11][9] ), .B2(n2823), .ZN(n1353) );
  OAI221_X1 U1250 ( .B1(n2880), .B2(n1301), .C1(n2877), .C2(n1302), .A(n1303), 
        .ZN(n1296) );
  AOI22_X1 U1251 ( .A1(\REGISTERS[26][10] ), .A2(n2874), .B1(
        \REGISTERS[27][10] ), .B2(n2871), .ZN(n1303) );
  OAI221_X1 U1252 ( .B1(n2832), .B2(n1317), .C1(n2829), .C2(n1318), .A(n1319), 
        .ZN(n1312) );
  AOI22_X1 U1253 ( .A1(\REGISTERS[10][10] ), .A2(n2826), .B1(
        \REGISTERS[11][10] ), .B2(n2823), .ZN(n1319) );
  OAI221_X1 U1254 ( .B1(n2880), .B2(n1267), .C1(n2877), .C2(n1268), .A(n1269), 
        .ZN(n1262) );
  AOI22_X1 U1255 ( .A1(\REGISTERS[26][11] ), .A2(n2874), .B1(
        \REGISTERS[27][11] ), .B2(n2871), .ZN(n1269) );
  OAI221_X1 U1256 ( .B1(n2832), .B2(n1283), .C1(n2829), .C2(n1284), .A(n1285), 
        .ZN(n1278) );
  AOI22_X1 U1257 ( .A1(\REGISTERS[10][11] ), .A2(n2826), .B1(
        \REGISTERS[11][11] ), .B2(n2823), .ZN(n1285) );
  OAI221_X1 U1258 ( .B1(n2881), .B2(n1233), .C1(n2878), .C2(n1234), .A(n1235), 
        .ZN(n1228) );
  AOI22_X1 U1259 ( .A1(\REGISTERS[26][12] ), .A2(n2875), .B1(
        \REGISTERS[27][12] ), .B2(n2872), .ZN(n1235) );
  OAI221_X1 U1260 ( .B1(n2833), .B2(n1249), .C1(n2830), .C2(n1250), .A(n1251), 
        .ZN(n1244) );
  AOI22_X1 U1261 ( .A1(\REGISTERS[10][12] ), .A2(n2827), .B1(
        \REGISTERS[11][12] ), .B2(n2824), .ZN(n1251) );
  OAI221_X1 U1262 ( .B1(n2881), .B2(n1199), .C1(n2878), .C2(n1200), .A(n1201), 
        .ZN(n1194) );
  AOI22_X1 U1263 ( .A1(\REGISTERS[26][13] ), .A2(n2875), .B1(
        \REGISTERS[27][13] ), .B2(n2872), .ZN(n1201) );
  OAI221_X1 U1264 ( .B1(n2833), .B2(n1215), .C1(n2830), .C2(n1216), .A(n1217), 
        .ZN(n1210) );
  AOI22_X1 U1265 ( .A1(\REGISTERS[10][13] ), .A2(n2827), .B1(
        \REGISTERS[11][13] ), .B2(n2824), .ZN(n1217) );
  OAI221_X1 U1266 ( .B1(n2881), .B2(n1165), .C1(n2878), .C2(n1166), .A(n1167), 
        .ZN(n1160) );
  AOI22_X1 U1267 ( .A1(\REGISTERS[26][14] ), .A2(n2875), .B1(
        \REGISTERS[27][14] ), .B2(n2872), .ZN(n1167) );
  OAI221_X1 U1268 ( .B1(n2833), .B2(n1181), .C1(n2830), .C2(n1182), .A(n1183), 
        .ZN(n1176) );
  AOI22_X1 U1269 ( .A1(\REGISTERS[10][14] ), .A2(n2827), .B1(
        \REGISTERS[11][14] ), .B2(n2824), .ZN(n1183) );
  OAI221_X1 U1270 ( .B1(n2881), .B2(n1131), .C1(n2878), .C2(n1132), .A(n1133), 
        .ZN(n1126) );
  AOI22_X1 U1271 ( .A1(\REGISTERS[26][15] ), .A2(n2875), .B1(
        \REGISTERS[27][15] ), .B2(n2872), .ZN(n1133) );
  OAI221_X1 U1272 ( .B1(n2833), .B2(n1147), .C1(n2830), .C2(n1148), .A(n1149), 
        .ZN(n1142) );
  AOI22_X1 U1273 ( .A1(\REGISTERS[10][15] ), .A2(n2827), .B1(
        \REGISTERS[11][15] ), .B2(n2824), .ZN(n1149) );
  OAI221_X1 U1274 ( .B1(n2881), .B2(n1097), .C1(n2878), .C2(n1098), .A(n1099), 
        .ZN(n1092) );
  AOI22_X1 U1275 ( .A1(\REGISTERS[26][16] ), .A2(n2875), .B1(
        \REGISTERS[27][16] ), .B2(n2872), .ZN(n1099) );
  OAI221_X1 U1276 ( .B1(n2833), .B2(n1113), .C1(n2830), .C2(n1114), .A(n1115), 
        .ZN(n1108) );
  AOI22_X1 U1277 ( .A1(\REGISTERS[10][16] ), .A2(n2827), .B1(
        \REGISTERS[11][16] ), .B2(n2824), .ZN(n1115) );
  OAI221_X1 U1278 ( .B1(n2881), .B2(n1063), .C1(n2878), .C2(n1064), .A(n1065), 
        .ZN(n1058) );
  AOI22_X1 U1279 ( .A1(\REGISTERS[26][17] ), .A2(n2875), .B1(
        \REGISTERS[27][17] ), .B2(n2872), .ZN(n1065) );
  OAI221_X1 U1280 ( .B1(n2833), .B2(n1079), .C1(n2830), .C2(n1080), .A(n1081), 
        .ZN(n1074) );
  AOI22_X1 U1281 ( .A1(\REGISTERS[10][17] ), .A2(n2827), .B1(
        \REGISTERS[11][17] ), .B2(n2824), .ZN(n1081) );
  OAI221_X1 U1282 ( .B1(n2881), .B2(n1029), .C1(n2878), .C2(n1030), .A(n1031), 
        .ZN(n1024) );
  AOI22_X1 U1283 ( .A1(\REGISTERS[26][18] ), .A2(n2875), .B1(
        \REGISTERS[27][18] ), .B2(n2872), .ZN(n1031) );
  OAI221_X1 U1284 ( .B1(n2833), .B2(n1045), .C1(n2830), .C2(n1046), .A(n1047), 
        .ZN(n1040) );
  AOI22_X1 U1285 ( .A1(\REGISTERS[10][18] ), .A2(n2827), .B1(
        \REGISTERS[11][18] ), .B2(n2824), .ZN(n1047) );
  OAI221_X1 U1286 ( .B1(n2881), .B2(n995), .C1(n2878), .C2(n996), .A(n997), 
        .ZN(n990) );
  AOI22_X1 U1287 ( .A1(\REGISTERS[26][19] ), .A2(n2875), .B1(
        \REGISTERS[27][19] ), .B2(n2872), .ZN(n997) );
  OAI221_X1 U1288 ( .B1(n2833), .B2(n1011), .C1(n2830), .C2(n1012), .A(n1013), 
        .ZN(n1006) );
  AOI22_X1 U1289 ( .A1(\REGISTERS[10][19] ), .A2(n2827), .B1(
        \REGISTERS[11][19] ), .B2(n2824), .ZN(n1013) );
  OAI221_X1 U1290 ( .B1(n2881), .B2(n961), .C1(n2878), .C2(n962), .A(n963), 
        .ZN(n956) );
  AOI22_X1 U1291 ( .A1(\REGISTERS[26][20] ), .A2(n2875), .B1(
        \REGISTERS[27][20] ), .B2(n2872), .ZN(n963) );
  OAI221_X1 U1292 ( .B1(n2833), .B2(n977), .C1(n2830), .C2(n978), .A(n979), 
        .ZN(n972) );
  AOI22_X1 U1293 ( .A1(\REGISTERS[10][20] ), .A2(n2827), .B1(
        \REGISTERS[11][20] ), .B2(n2824), .ZN(n979) );
  OAI221_X1 U1294 ( .B1(n2881), .B2(n927), .C1(n2878), .C2(n928), .A(n929), 
        .ZN(n922) );
  AOI22_X1 U1295 ( .A1(\REGISTERS[26][21] ), .A2(n2875), .B1(
        \REGISTERS[27][21] ), .B2(n2872), .ZN(n929) );
  OAI221_X1 U1296 ( .B1(n2833), .B2(n943), .C1(n2830), .C2(n944), .A(n945), 
        .ZN(n938) );
  AOI22_X1 U1297 ( .A1(\REGISTERS[10][21] ), .A2(n2827), .B1(
        \REGISTERS[11][21] ), .B2(n2824), .ZN(n945) );
  OAI221_X1 U1298 ( .B1(n2881), .B2(n893), .C1(n2878), .C2(n894), .A(n895), 
        .ZN(n888) );
  AOI22_X1 U1299 ( .A1(\REGISTERS[26][22] ), .A2(n2875), .B1(
        \REGISTERS[27][22] ), .B2(n2872), .ZN(n895) );
  OAI221_X1 U1300 ( .B1(n2833), .B2(n909), .C1(n2830), .C2(n910), .A(n911), 
        .ZN(n904) );
  AOI22_X1 U1301 ( .A1(\REGISTERS[10][22] ), .A2(n2827), .B1(
        \REGISTERS[11][22] ), .B2(n2824), .ZN(n911) );
  OAI221_X1 U1302 ( .B1(n2881), .B2(n859), .C1(n2878), .C2(n860), .A(n861), 
        .ZN(n854) );
  AOI22_X1 U1303 ( .A1(\REGISTERS[26][23] ), .A2(n2875), .B1(
        \REGISTERS[27][23] ), .B2(n2872), .ZN(n861) );
  OAI221_X1 U1304 ( .B1(n2833), .B2(n875), .C1(n2830), .C2(n876), .A(n877), 
        .ZN(n870) );
  AOI22_X1 U1305 ( .A1(\REGISTERS[10][23] ), .A2(n2827), .B1(
        \REGISTERS[11][23] ), .B2(n2824), .ZN(n877) );
  OAI221_X1 U1306 ( .B1(n2870), .B2(n828), .C1(n2867), .C2(n829), .A(n830), 
        .ZN(n819) );
  AOI22_X1 U1307 ( .A1(\REGISTERS[22][24] ), .A2(n2864), .B1(
        \REGISTERS[23][24] ), .B2(n2861), .ZN(n830) );
  OAI221_X1 U1308 ( .B1(n2822), .B2(n844), .C1(n2819), .C2(n845), .A(n846), 
        .ZN(n835) );
  AOI22_X1 U1309 ( .A1(\REGISTERS[6][24] ), .A2(n2816), .B1(\REGISTERS[7][24] ), .B2(n2813), .ZN(n846) );
  OAI221_X1 U1310 ( .B1(n2870), .B2(n794), .C1(n2867), .C2(n795), .A(n796), 
        .ZN(n785) );
  AOI22_X1 U1311 ( .A1(\REGISTERS[22][25] ), .A2(n2864), .B1(
        \REGISTERS[23][25] ), .B2(n2861), .ZN(n796) );
  OAI221_X1 U1312 ( .B1(n2822), .B2(n810), .C1(n2819), .C2(n811), .A(n812), 
        .ZN(n801) );
  AOI22_X1 U1313 ( .A1(\REGISTERS[6][25] ), .A2(n2816), .B1(\REGISTERS[7][25] ), .B2(n2813), .ZN(n812) );
  OAI221_X1 U1314 ( .B1(n2870), .B2(n760), .C1(n2867), .C2(n761), .A(n762), 
        .ZN(n751) );
  AOI22_X1 U1315 ( .A1(\REGISTERS[22][26] ), .A2(n2864), .B1(
        \REGISTERS[23][26] ), .B2(n2861), .ZN(n762) );
  OAI221_X1 U1316 ( .B1(n2822), .B2(n776), .C1(n2819), .C2(n777), .A(n778), 
        .ZN(n767) );
  AOI22_X1 U1317 ( .A1(\REGISTERS[6][26] ), .A2(n2816), .B1(\REGISTERS[7][26] ), .B2(n2813), .ZN(n778) );
  OAI221_X1 U1318 ( .B1(n2870), .B2(n726), .C1(n2867), .C2(n727), .A(n728), 
        .ZN(n717) );
  AOI22_X1 U1319 ( .A1(\REGISTERS[22][27] ), .A2(n2864), .B1(
        \REGISTERS[23][27] ), .B2(n2861), .ZN(n728) );
  OAI221_X1 U1320 ( .B1(n2822), .B2(n742), .C1(n2819), .C2(n743), .A(n744), 
        .ZN(n733) );
  AOI22_X1 U1321 ( .A1(\REGISTERS[6][27] ), .A2(n2816), .B1(\REGISTERS[7][27] ), .B2(n2813), .ZN(n744) );
  OAI221_X1 U1322 ( .B1(n2870), .B2(n692), .C1(n2867), .C2(n693), .A(n694), 
        .ZN(n683) );
  AOI22_X1 U1323 ( .A1(\REGISTERS[22][28] ), .A2(n2864), .B1(
        \REGISTERS[23][28] ), .B2(n2861), .ZN(n694) );
  OAI221_X1 U1324 ( .B1(n2822), .B2(n708), .C1(n2819), .C2(n709), .A(n710), 
        .ZN(n699) );
  AOI22_X1 U1325 ( .A1(\REGISTERS[6][28] ), .A2(n2816), .B1(\REGISTERS[7][28] ), .B2(n2813), .ZN(n710) );
  OAI221_X1 U1326 ( .B1(n2870), .B2(n658), .C1(n2867), .C2(n659), .A(n660), 
        .ZN(n649) );
  AOI22_X1 U1327 ( .A1(\REGISTERS[22][29] ), .A2(n2864), .B1(
        \REGISTERS[23][29] ), .B2(n2861), .ZN(n660) );
  OAI221_X1 U1328 ( .B1(n2822), .B2(n674), .C1(n2819), .C2(n675), .A(n676), 
        .ZN(n665) );
  AOI22_X1 U1329 ( .A1(\REGISTERS[6][29] ), .A2(n2816), .B1(\REGISTERS[7][29] ), .B2(n2813), .ZN(n676) );
  OAI221_X1 U1330 ( .B1(n2870), .B2(n624), .C1(n2867), .C2(n625), .A(n626), 
        .ZN(n615) );
  AOI22_X1 U1331 ( .A1(\REGISTERS[22][30] ), .A2(n2864), .B1(
        \REGISTERS[23][30] ), .B2(n2861), .ZN(n626) );
  OAI221_X1 U1332 ( .B1(n2822), .B2(n640), .C1(n2819), .C2(n641), .A(n642), 
        .ZN(n631) );
  AOI22_X1 U1333 ( .A1(\REGISTERS[6][30] ), .A2(n2816), .B1(\REGISTERS[7][30] ), .B2(n2813), .ZN(n642) );
  OAI221_X1 U1334 ( .B1(n2870), .B2(n567), .C1(n2867), .C2(n569), .A(n570), 
        .ZN(n549) );
  AOI22_X1 U1335 ( .A1(\REGISTERS[22][31] ), .A2(n2864), .B1(
        \REGISTERS[23][31] ), .B2(n2861), .ZN(n570) );
  OAI221_X1 U1336 ( .B1(n2822), .B2(n599), .C1(n2819), .C2(n601), .A(n602), 
        .ZN(n581) );
  AOI22_X1 U1337 ( .A1(\REGISTERS[6][31] ), .A2(n2816), .B1(\REGISTERS[7][31] ), .B2(n2813), .ZN(n602) );
  OAI221_X1 U1338 ( .B1(n2858), .B2(n831), .C1(n2855), .C2(n832), .A(n833), 
        .ZN(n818) );
  AOI22_X1 U1339 ( .A1(\REGISTERS[18][24] ), .A2(n2852), .B1(
        \REGISTERS[19][24] ), .B2(n2849), .ZN(n833) );
  OAI221_X1 U1340 ( .B1(n2858), .B2(n797), .C1(n2855), .C2(n798), .A(n799), 
        .ZN(n784) );
  AOI22_X1 U1341 ( .A1(\REGISTERS[18][25] ), .A2(n2852), .B1(
        \REGISTERS[19][25] ), .B2(n2849), .ZN(n799) );
  OAI221_X1 U1342 ( .B1(n2858), .B2(n763), .C1(n2855), .C2(n764), .A(n765), 
        .ZN(n750) );
  AOI22_X1 U1343 ( .A1(\REGISTERS[18][26] ), .A2(n2852), .B1(
        \REGISTERS[19][26] ), .B2(n2849), .ZN(n765) );
  OAI221_X1 U1344 ( .B1(n2858), .B2(n729), .C1(n2855), .C2(n730), .A(n731), 
        .ZN(n716) );
  AOI22_X1 U1345 ( .A1(\REGISTERS[18][27] ), .A2(n2852), .B1(
        \REGISTERS[19][27] ), .B2(n2849), .ZN(n731) );
  OAI221_X1 U1346 ( .B1(n2858), .B2(n695), .C1(n2855), .C2(n696), .A(n697), 
        .ZN(n682) );
  AOI22_X1 U1347 ( .A1(\REGISTERS[18][28] ), .A2(n2852), .B1(
        \REGISTERS[19][28] ), .B2(n2849), .ZN(n697) );
  OAI221_X1 U1348 ( .B1(n2858), .B2(n661), .C1(n2855), .C2(n662), .A(n663), 
        .ZN(n648) );
  AOI22_X1 U1349 ( .A1(\REGISTERS[18][29] ), .A2(n2852), .B1(
        \REGISTERS[19][29] ), .B2(n2849), .ZN(n663) );
  OAI221_X1 U1350 ( .B1(n2858), .B2(n627), .C1(n2855), .C2(n628), .A(n629), 
        .ZN(n614) );
  AOI22_X1 U1351 ( .A1(\REGISTERS[18][30] ), .A2(n2852), .B1(
        \REGISTERS[19][30] ), .B2(n2849), .ZN(n629) );
  OAI221_X1 U1352 ( .B1(n2858), .B2(n574), .C1(n2855), .C2(n576), .A(n577), 
        .ZN(n548) );
  AOI22_X1 U1353 ( .A1(\REGISTERS[18][31] ), .A2(n2852), .B1(
        \REGISTERS[19][31] ), .B2(n2849), .ZN(n577) );
  OAI221_X1 U1354 ( .B1(n828), .B2(n2774), .C1(n829), .C2(n2771), .A(n1848), 
        .ZN(n1843) );
  AOI22_X1 U1355 ( .A1(n2768), .A2(\REGISTERS[22][24] ), .B1(n2763), .B2(
        \REGISTERS[23][24] ), .ZN(n1848) );
  OAI221_X1 U1356 ( .B1(n844), .B2(n2726), .C1(n845), .C2(n2723), .A(n1856), 
        .ZN(n1851) );
  AOI22_X1 U1357 ( .A1(n2720), .A2(\REGISTERS[6][24] ), .B1(n2715), .B2(
        \REGISTERS[7][24] ), .ZN(n1856) );
  OAI221_X1 U1358 ( .B1(n794), .B2(n2774), .C1(n795), .C2(n2771), .A(n1830), 
        .ZN(n1825) );
  AOI22_X1 U1359 ( .A1(n2768), .A2(\REGISTERS[22][25] ), .B1(n2763), .B2(
        \REGISTERS[23][25] ), .ZN(n1830) );
  OAI221_X1 U1360 ( .B1(n810), .B2(n2726), .C1(n811), .C2(n2723), .A(n1838), 
        .ZN(n1833) );
  AOI22_X1 U1361 ( .A1(n2720), .A2(\REGISTERS[6][25] ), .B1(n2715), .B2(
        \REGISTERS[7][25] ), .ZN(n1838) );
  OAI221_X1 U1362 ( .B1(n760), .B2(n2774), .C1(n761), .C2(n2771), .A(n1812), 
        .ZN(n1807) );
  AOI22_X1 U1363 ( .A1(n2768), .A2(\REGISTERS[22][26] ), .B1(n2763), .B2(
        \REGISTERS[23][26] ), .ZN(n1812) );
  OAI221_X1 U1364 ( .B1(n776), .B2(n2726), .C1(n777), .C2(n2723), .A(n1820), 
        .ZN(n1815) );
  AOI22_X1 U1365 ( .A1(n2720), .A2(\REGISTERS[6][26] ), .B1(n2715), .B2(
        \REGISTERS[7][26] ), .ZN(n1820) );
  OAI221_X1 U1366 ( .B1(n726), .B2(n2774), .C1(n727), .C2(n2771), .A(n1794), 
        .ZN(n1789) );
  AOI22_X1 U1367 ( .A1(n2768), .A2(\REGISTERS[22][27] ), .B1(n2763), .B2(
        \REGISTERS[23][27] ), .ZN(n1794) );
  OAI221_X1 U1368 ( .B1(n742), .B2(n2726), .C1(n743), .C2(n2723), .A(n1802), 
        .ZN(n1797) );
  AOI22_X1 U1369 ( .A1(n2720), .A2(\REGISTERS[6][27] ), .B1(n2715), .B2(
        \REGISTERS[7][27] ), .ZN(n1802) );
  OAI221_X1 U1370 ( .B1(n692), .B2(n2774), .C1(n693), .C2(n2771), .A(n1776), 
        .ZN(n1771) );
  AOI22_X1 U1371 ( .A1(n2768), .A2(\REGISTERS[22][28] ), .B1(n2763), .B2(
        \REGISTERS[23][28] ), .ZN(n1776) );
  OAI221_X1 U1372 ( .B1(n708), .B2(n2726), .C1(n709), .C2(n2723), .A(n1784), 
        .ZN(n1779) );
  AOI22_X1 U1373 ( .A1(n2720), .A2(\REGISTERS[6][28] ), .B1(n2715), .B2(
        \REGISTERS[7][28] ), .ZN(n1784) );
  OAI221_X1 U1374 ( .B1(n658), .B2(n2774), .C1(n659), .C2(n2771), .A(n1758), 
        .ZN(n1753) );
  AOI22_X1 U1375 ( .A1(n2768), .A2(\REGISTERS[22][29] ), .B1(n2763), .B2(
        \REGISTERS[23][29] ), .ZN(n1758) );
  OAI221_X1 U1376 ( .B1(n674), .B2(n2726), .C1(n675), .C2(n2723), .A(n1766), 
        .ZN(n1761) );
  AOI22_X1 U1377 ( .A1(n2720), .A2(\REGISTERS[6][29] ), .B1(n2715), .B2(
        \REGISTERS[7][29] ), .ZN(n1766) );
  OAI221_X1 U1378 ( .B1(n624), .B2(n2774), .C1(n625), .C2(n2771), .A(n1740), 
        .ZN(n1735) );
  AOI22_X1 U1379 ( .A1(n2768), .A2(\REGISTERS[22][30] ), .B1(n2763), .B2(
        \REGISTERS[23][30] ), .ZN(n1740) );
  OAI221_X1 U1380 ( .B1(n640), .B2(n2726), .C1(n641), .C2(n2723), .A(n1748), 
        .ZN(n1743) );
  AOI22_X1 U1381 ( .A1(n2720), .A2(\REGISTERS[6][30] ), .B1(n2715), .B2(
        \REGISTERS[7][30] ), .ZN(n1748) );
  OAI221_X1 U1382 ( .B1(n567), .B2(n2774), .C1(n569), .C2(n2771), .A(n1700), 
        .ZN(n1685) );
  AOI22_X1 U1383 ( .A1(n2768), .A2(\REGISTERS[22][31] ), .B1(n2763), .B2(
        \REGISTERS[23][31] ), .ZN(n1700) );
  OAI221_X1 U1384 ( .B1(n599), .B2(n2726), .C1(n601), .C2(n2723), .A(n1724), 
        .ZN(n1709) );
  AOI22_X1 U1385 ( .A1(n2720), .A2(\REGISTERS[6][31] ), .B1(n2715), .B2(
        \REGISTERS[7][31] ), .ZN(n1724) );
  OAI221_X1 U1386 ( .B1(n831), .B2(n2762), .C1(n832), .C2(n2759), .A(n1849), 
        .ZN(n1842) );
  AOI22_X1 U1387 ( .A1(n2756), .A2(\REGISTERS[18][24] ), .B1(n2751), .B2(
        \REGISTERS[19][24] ), .ZN(n1849) );
  OAI221_X1 U1388 ( .B1(n797), .B2(n2762), .C1(n798), .C2(n2759), .A(n1831), 
        .ZN(n1824) );
  AOI22_X1 U1389 ( .A1(n2756), .A2(\REGISTERS[18][25] ), .B1(n2751), .B2(
        \REGISTERS[19][25] ), .ZN(n1831) );
  OAI221_X1 U1390 ( .B1(n763), .B2(n2762), .C1(n764), .C2(n2759), .A(n1813), 
        .ZN(n1806) );
  AOI22_X1 U1391 ( .A1(n2756), .A2(\REGISTERS[18][26] ), .B1(n2751), .B2(
        \REGISTERS[19][26] ), .ZN(n1813) );
  OAI221_X1 U1392 ( .B1(n729), .B2(n2762), .C1(n730), .C2(n2759), .A(n1795), 
        .ZN(n1788) );
  AOI22_X1 U1393 ( .A1(n2756), .A2(\REGISTERS[18][27] ), .B1(n2751), .B2(
        \REGISTERS[19][27] ), .ZN(n1795) );
  OAI221_X1 U1394 ( .B1(n695), .B2(n2762), .C1(n696), .C2(n2759), .A(n1777), 
        .ZN(n1770) );
  AOI22_X1 U1395 ( .A1(n2756), .A2(\REGISTERS[18][28] ), .B1(n2751), .B2(
        \REGISTERS[19][28] ), .ZN(n1777) );
  OAI221_X1 U1396 ( .B1(n661), .B2(n2762), .C1(n662), .C2(n2759), .A(n1759), 
        .ZN(n1752) );
  AOI22_X1 U1397 ( .A1(n2756), .A2(\REGISTERS[18][29] ), .B1(n2751), .B2(
        \REGISTERS[19][29] ), .ZN(n1759) );
  OAI221_X1 U1398 ( .B1(n627), .B2(n2762), .C1(n628), .C2(n2759), .A(n1741), 
        .ZN(n1734) );
  AOI22_X1 U1399 ( .A1(n2756), .A2(\REGISTERS[18][30] ), .B1(n2751), .B2(
        \REGISTERS[19][30] ), .ZN(n1741) );
  OAI221_X1 U1400 ( .B1(n574), .B2(n2762), .C1(n576), .C2(n2759), .A(n1705), 
        .ZN(n1684) );
  AOI22_X1 U1401 ( .A1(n2756), .A2(\REGISTERS[18][31] ), .B1(n2751), .B2(
        \REGISTERS[19][31] ), .ZN(n1705) );
  OAI221_X1 U1402 ( .B1(n1651), .B2(n2772), .C1(n1652), .C2(n2769), .A(n2287), 
        .ZN(n2275) );
  AOI22_X1 U1403 ( .A1(n2766), .A2(\REGISTERS[22][0] ), .B1(n2765), .B2(
        \REGISTERS[23][0] ), .ZN(n2287) );
  OAI221_X1 U1404 ( .B1(n1672), .B2(n2724), .C1(n1673), .C2(n2721), .A(n2300), 
        .ZN(n2293) );
  AOI22_X1 U1405 ( .A1(n2718), .A2(\REGISTERS[6][0] ), .B1(n2717), .B2(
        \REGISTERS[7][0] ), .ZN(n2300) );
  OAI221_X1 U1406 ( .B1(n1610), .B2(n2772), .C1(n1611), .C2(n2769), .A(n2262), 
        .ZN(n2257) );
  AOI22_X1 U1407 ( .A1(n2766), .A2(\REGISTERS[22][1] ), .B1(n2765), .B2(
        \REGISTERS[23][1] ), .ZN(n2262) );
  OAI221_X1 U1408 ( .B1(n1626), .B2(n2724), .C1(n1627), .C2(n2721), .A(n2270), 
        .ZN(n2265) );
  AOI22_X1 U1409 ( .A1(n2718), .A2(\REGISTERS[6][1] ), .B1(n2717), .B2(
        \REGISTERS[7][1] ), .ZN(n2270) );
  OAI221_X1 U1410 ( .B1(n1576), .B2(n2772), .C1(n1577), .C2(n2769), .A(n2244), 
        .ZN(n2239) );
  AOI22_X1 U1411 ( .A1(n2766), .A2(\REGISTERS[22][2] ), .B1(n2765), .B2(
        \REGISTERS[23][2] ), .ZN(n2244) );
  OAI221_X1 U1412 ( .B1(n1592), .B2(n2724), .C1(n1593), .C2(n2721), .A(n2252), 
        .ZN(n2247) );
  AOI22_X1 U1413 ( .A1(n2718), .A2(\REGISTERS[6][2] ), .B1(n2717), .B2(
        \REGISTERS[7][2] ), .ZN(n2252) );
  OAI221_X1 U1414 ( .B1(n1542), .B2(n2772), .C1(n1543), .C2(n2769), .A(n2226), 
        .ZN(n2221) );
  AOI22_X1 U1415 ( .A1(n2766), .A2(\REGISTERS[22][3] ), .B1(n2765), .B2(
        \REGISTERS[23][3] ), .ZN(n2226) );
  OAI221_X1 U1416 ( .B1(n1558), .B2(n2724), .C1(n1559), .C2(n2721), .A(n2234), 
        .ZN(n2229) );
  AOI22_X1 U1417 ( .A1(n2718), .A2(\REGISTERS[6][3] ), .B1(n2717), .B2(
        \REGISTERS[7][3] ), .ZN(n2234) );
  OAI221_X1 U1418 ( .B1(n1508), .B2(n2772), .C1(n1509), .C2(n2769), .A(n2208), 
        .ZN(n2203) );
  AOI22_X1 U1419 ( .A1(n2766), .A2(\REGISTERS[22][4] ), .B1(n2765), .B2(
        \REGISTERS[23][4] ), .ZN(n2208) );
  OAI221_X1 U1420 ( .B1(n1524), .B2(n2724), .C1(n1525), .C2(n2721), .A(n2216), 
        .ZN(n2211) );
  AOI22_X1 U1421 ( .A1(n2718), .A2(\REGISTERS[6][4] ), .B1(n2717), .B2(
        \REGISTERS[7][4] ), .ZN(n2216) );
  OAI221_X1 U1422 ( .B1(n1474), .B2(n2772), .C1(n1475), .C2(n2769), .A(n2190), 
        .ZN(n2185) );
  AOI22_X1 U1423 ( .A1(n2766), .A2(\REGISTERS[22][5] ), .B1(n2765), .B2(
        \REGISTERS[23][5] ), .ZN(n2190) );
  OAI221_X1 U1424 ( .B1(n1490), .B2(n2724), .C1(n1491), .C2(n2721), .A(n2198), 
        .ZN(n2193) );
  AOI22_X1 U1425 ( .A1(n2718), .A2(\REGISTERS[6][5] ), .B1(n2717), .B2(
        \REGISTERS[7][5] ), .ZN(n2198) );
  OAI221_X1 U1426 ( .B1(n1440), .B2(n2772), .C1(n1441), .C2(n2769), .A(n2172), 
        .ZN(n2167) );
  AOI22_X1 U1427 ( .A1(n2766), .A2(\REGISTERS[22][6] ), .B1(n2765), .B2(
        \REGISTERS[23][6] ), .ZN(n2172) );
  OAI221_X1 U1428 ( .B1(n1456), .B2(n2724), .C1(n1457), .C2(n2721), .A(n2180), 
        .ZN(n2175) );
  AOI22_X1 U1429 ( .A1(n2718), .A2(\REGISTERS[6][6] ), .B1(n2717), .B2(
        \REGISTERS[7][6] ), .ZN(n2180) );
  OAI221_X1 U1430 ( .B1(n1406), .B2(n2772), .C1(n1407), .C2(n2769), .A(n2154), 
        .ZN(n2149) );
  AOI22_X1 U1431 ( .A1(n2766), .A2(\REGISTERS[22][7] ), .B1(n2765), .B2(
        \REGISTERS[23][7] ), .ZN(n2154) );
  OAI221_X1 U1432 ( .B1(n1422), .B2(n2724), .C1(n1423), .C2(n2721), .A(n2162), 
        .ZN(n2157) );
  AOI22_X1 U1433 ( .A1(n2718), .A2(\REGISTERS[6][7] ), .B1(n2717), .B2(
        \REGISTERS[7][7] ), .ZN(n2162) );
  OAI221_X1 U1434 ( .B1(n1372), .B2(n2772), .C1(n1373), .C2(n2769), .A(n2136), 
        .ZN(n2131) );
  AOI22_X1 U1435 ( .A1(n2766), .A2(\REGISTERS[22][8] ), .B1(n2764), .B2(
        \REGISTERS[23][8] ), .ZN(n2136) );
  OAI221_X1 U1436 ( .B1(n1388), .B2(n2724), .C1(n1389), .C2(n2721), .A(n2144), 
        .ZN(n2139) );
  AOI22_X1 U1437 ( .A1(n2718), .A2(\REGISTERS[6][8] ), .B1(n2716), .B2(
        \REGISTERS[7][8] ), .ZN(n2144) );
  OAI221_X1 U1438 ( .B1(n1338), .B2(n2772), .C1(n1339), .C2(n2769), .A(n2118), 
        .ZN(n2113) );
  AOI22_X1 U1439 ( .A1(n2766), .A2(\REGISTERS[22][9] ), .B1(n2764), .B2(
        \REGISTERS[23][9] ), .ZN(n2118) );
  OAI221_X1 U1440 ( .B1(n1354), .B2(n2724), .C1(n1355), .C2(n2721), .A(n2126), 
        .ZN(n2121) );
  AOI22_X1 U1441 ( .A1(n2718), .A2(\REGISTERS[6][9] ), .B1(n2716), .B2(
        \REGISTERS[7][9] ), .ZN(n2126) );
  OAI221_X1 U1442 ( .B1(n1304), .B2(n2772), .C1(n1305), .C2(n2769), .A(n2100), 
        .ZN(n2095) );
  AOI22_X1 U1443 ( .A1(n2766), .A2(\REGISTERS[22][10] ), .B1(n2764), .B2(
        \REGISTERS[23][10] ), .ZN(n2100) );
  OAI221_X1 U1444 ( .B1(n1320), .B2(n2724), .C1(n1321), .C2(n2721), .A(n2108), 
        .ZN(n2103) );
  AOI22_X1 U1445 ( .A1(n2718), .A2(\REGISTERS[6][10] ), .B1(n2716), .B2(
        \REGISTERS[7][10] ), .ZN(n2108) );
  OAI221_X1 U1446 ( .B1(n1270), .B2(n2772), .C1(n1271), .C2(n2769), .A(n2082), 
        .ZN(n2077) );
  AOI22_X1 U1447 ( .A1(n2766), .A2(\REGISTERS[22][11] ), .B1(n2764), .B2(
        \REGISTERS[23][11] ), .ZN(n2082) );
  OAI221_X1 U1448 ( .B1(n1286), .B2(n2724), .C1(n1287), .C2(n2721), .A(n2090), 
        .ZN(n2085) );
  AOI22_X1 U1449 ( .A1(n2718), .A2(\REGISTERS[6][11] ), .B1(n2716), .B2(
        \REGISTERS[7][11] ), .ZN(n2090) );
  OAI221_X1 U1450 ( .B1(n1236), .B2(n2773), .C1(n1237), .C2(n2770), .A(n2064), 
        .ZN(n2059) );
  AOI22_X1 U1451 ( .A1(n2767), .A2(\REGISTERS[22][12] ), .B1(n2764), .B2(
        \REGISTERS[23][12] ), .ZN(n2064) );
  OAI221_X1 U1452 ( .B1(n1252), .B2(n2725), .C1(n1253), .C2(n2722), .A(n2072), 
        .ZN(n2067) );
  AOI22_X1 U1453 ( .A1(n2719), .A2(\REGISTERS[6][12] ), .B1(n2716), .B2(
        \REGISTERS[7][12] ), .ZN(n2072) );
  OAI221_X1 U1454 ( .B1(n1202), .B2(n2773), .C1(n1203), .C2(n2770), .A(n2046), 
        .ZN(n2041) );
  AOI22_X1 U1455 ( .A1(n2767), .A2(\REGISTERS[22][13] ), .B1(n2764), .B2(
        \REGISTERS[23][13] ), .ZN(n2046) );
  OAI221_X1 U1456 ( .B1(n1218), .B2(n2725), .C1(n1219), .C2(n2722), .A(n2054), 
        .ZN(n2049) );
  AOI22_X1 U1457 ( .A1(n2719), .A2(\REGISTERS[6][13] ), .B1(n2716), .B2(
        \REGISTERS[7][13] ), .ZN(n2054) );
  OAI221_X1 U1458 ( .B1(n1168), .B2(n2773), .C1(n1169), .C2(n2770), .A(n2028), 
        .ZN(n2023) );
  AOI22_X1 U1459 ( .A1(n2767), .A2(\REGISTERS[22][14] ), .B1(n2764), .B2(
        \REGISTERS[23][14] ), .ZN(n2028) );
  OAI221_X1 U1460 ( .B1(n1184), .B2(n2725), .C1(n1185), .C2(n2722), .A(n2036), 
        .ZN(n2031) );
  AOI22_X1 U1461 ( .A1(n2719), .A2(\REGISTERS[6][14] ), .B1(n2716), .B2(
        \REGISTERS[7][14] ), .ZN(n2036) );
  OAI221_X1 U1462 ( .B1(n1134), .B2(n2773), .C1(n1135), .C2(n2770), .A(n2010), 
        .ZN(n2005) );
  AOI22_X1 U1463 ( .A1(n2767), .A2(\REGISTERS[22][15] ), .B1(n2764), .B2(
        \REGISTERS[23][15] ), .ZN(n2010) );
  OAI221_X1 U1464 ( .B1(n1150), .B2(n2725), .C1(n1151), .C2(n2722), .A(n2018), 
        .ZN(n2013) );
  AOI22_X1 U1465 ( .A1(n2719), .A2(\REGISTERS[6][15] ), .B1(n2716), .B2(
        \REGISTERS[7][15] ), .ZN(n2018) );
  OAI221_X1 U1466 ( .B1(n1100), .B2(n2773), .C1(n1101), .C2(n2770), .A(n1992), 
        .ZN(n1987) );
  AOI22_X1 U1467 ( .A1(n2767), .A2(\REGISTERS[22][16] ), .B1(n2764), .B2(
        \REGISTERS[23][16] ), .ZN(n1992) );
  OAI221_X1 U1468 ( .B1(n1116), .B2(n2725), .C1(n1117), .C2(n2722), .A(n2000), 
        .ZN(n1995) );
  AOI22_X1 U1469 ( .A1(n2719), .A2(\REGISTERS[6][16] ), .B1(n2716), .B2(
        \REGISTERS[7][16] ), .ZN(n2000) );
  OAI221_X1 U1470 ( .B1(n1066), .B2(n2773), .C1(n1067), .C2(n2770), .A(n1974), 
        .ZN(n1969) );
  AOI22_X1 U1471 ( .A1(n2767), .A2(\REGISTERS[22][17] ), .B1(n2764), .B2(
        \REGISTERS[23][17] ), .ZN(n1974) );
  OAI221_X1 U1472 ( .B1(n1082), .B2(n2725), .C1(n1083), .C2(n2722), .A(n1982), 
        .ZN(n1977) );
  AOI22_X1 U1473 ( .A1(n2719), .A2(\REGISTERS[6][17] ), .B1(n2716), .B2(
        \REGISTERS[7][17] ), .ZN(n1982) );
  OAI221_X1 U1474 ( .B1(n1032), .B2(n2773), .C1(n1033), .C2(n2770), .A(n1956), 
        .ZN(n1951) );
  AOI22_X1 U1475 ( .A1(n2767), .A2(\REGISTERS[22][18] ), .B1(n2764), .B2(
        \REGISTERS[23][18] ), .ZN(n1956) );
  OAI221_X1 U1476 ( .B1(n1048), .B2(n2725), .C1(n1049), .C2(n2722), .A(n1964), 
        .ZN(n1959) );
  AOI22_X1 U1477 ( .A1(n2719), .A2(\REGISTERS[6][18] ), .B1(n2716), .B2(
        \REGISTERS[7][18] ), .ZN(n1964) );
  OAI221_X1 U1478 ( .B1(n998), .B2(n2773), .C1(n999), .C2(n2770), .A(n1938), 
        .ZN(n1933) );
  AOI22_X1 U1479 ( .A1(n2767), .A2(\REGISTERS[22][19] ), .B1(n2764), .B2(
        \REGISTERS[23][19] ), .ZN(n1938) );
  OAI221_X1 U1480 ( .B1(n1014), .B2(n2725), .C1(n1015), .C2(n2722), .A(n1946), 
        .ZN(n1941) );
  AOI22_X1 U1481 ( .A1(n2719), .A2(\REGISTERS[6][19] ), .B1(n2716), .B2(
        \REGISTERS[7][19] ), .ZN(n1946) );
  OAI221_X1 U1482 ( .B1(n964), .B2(n2773), .C1(n965), .C2(n2770), .A(n1920), 
        .ZN(n1915) );
  AOI22_X1 U1483 ( .A1(n2767), .A2(\REGISTERS[22][20] ), .B1(n2763), .B2(
        \REGISTERS[23][20] ), .ZN(n1920) );
  OAI221_X1 U1484 ( .B1(n980), .B2(n2725), .C1(n981), .C2(n2722), .A(n1928), 
        .ZN(n1923) );
  AOI22_X1 U1485 ( .A1(n2719), .A2(\REGISTERS[6][20] ), .B1(n2715), .B2(
        \REGISTERS[7][20] ), .ZN(n1928) );
  OAI221_X1 U1486 ( .B1(n930), .B2(n2773), .C1(n931), .C2(n2770), .A(n1902), 
        .ZN(n1897) );
  AOI22_X1 U1487 ( .A1(n2767), .A2(\REGISTERS[22][21] ), .B1(n2763), .B2(
        \REGISTERS[23][21] ), .ZN(n1902) );
  OAI221_X1 U1488 ( .B1(n946), .B2(n2725), .C1(n947), .C2(n2722), .A(n1910), 
        .ZN(n1905) );
  AOI22_X1 U1489 ( .A1(n2719), .A2(\REGISTERS[6][21] ), .B1(n2715), .B2(
        \REGISTERS[7][21] ), .ZN(n1910) );
  OAI221_X1 U1490 ( .B1(n896), .B2(n2773), .C1(n897), .C2(n2770), .A(n1884), 
        .ZN(n1879) );
  AOI22_X1 U1491 ( .A1(n2767), .A2(\REGISTERS[22][22] ), .B1(n2763), .B2(
        \REGISTERS[23][22] ), .ZN(n1884) );
  OAI221_X1 U1492 ( .B1(n912), .B2(n2725), .C1(n913), .C2(n2722), .A(n1892), 
        .ZN(n1887) );
  AOI22_X1 U1493 ( .A1(n2719), .A2(\REGISTERS[6][22] ), .B1(n2715), .B2(
        \REGISTERS[7][22] ), .ZN(n1892) );
  OAI221_X1 U1494 ( .B1(n862), .B2(n2773), .C1(n863), .C2(n2770), .A(n1866), 
        .ZN(n1861) );
  AOI22_X1 U1495 ( .A1(n2767), .A2(\REGISTERS[22][23] ), .B1(n2763), .B2(
        \REGISTERS[23][23] ), .ZN(n1866) );
  OAI221_X1 U1496 ( .B1(n878), .B2(n2725), .C1(n879), .C2(n2722), .A(n1874), 
        .ZN(n1869) );
  AOI22_X1 U1497 ( .A1(n2719), .A2(\REGISTERS[6][23] ), .B1(n2715), .B2(
        \REGISTERS[7][23] ), .ZN(n1874) );
  OAI221_X1 U1498 ( .B1(n2868), .B2(n1651), .C1(n2865), .C2(n1652), .A(n1653), 
        .ZN(n1635) );
  AOI22_X1 U1499 ( .A1(\REGISTERS[22][0] ), .A2(n2862), .B1(\REGISTERS[23][0] ), .B2(n2859), .ZN(n1653) );
  OAI221_X1 U1500 ( .B1(n2820), .B2(n1672), .C1(n2817), .C2(n1673), .A(n1674), 
        .ZN(n1661) );
  AOI22_X1 U1501 ( .A1(\REGISTERS[6][0] ), .A2(n2814), .B1(\REGISTERS[7][0] ), 
        .B2(n2811), .ZN(n1674) );
  OAI221_X1 U1502 ( .B1(n2868), .B2(n1610), .C1(n2865), .C2(n1611), .A(n1612), 
        .ZN(n1601) );
  AOI22_X1 U1503 ( .A1(\REGISTERS[22][1] ), .A2(n2862), .B1(\REGISTERS[23][1] ), .B2(n2859), .ZN(n1612) );
  OAI221_X1 U1504 ( .B1(n2820), .B2(n1626), .C1(n2817), .C2(n1627), .A(n1628), 
        .ZN(n1617) );
  AOI22_X1 U1505 ( .A1(\REGISTERS[6][1] ), .A2(n2814), .B1(\REGISTERS[7][1] ), 
        .B2(n2811), .ZN(n1628) );
  OAI221_X1 U1506 ( .B1(n2868), .B2(n1576), .C1(n2865), .C2(n1577), .A(n1578), 
        .ZN(n1567) );
  AOI22_X1 U1507 ( .A1(\REGISTERS[22][2] ), .A2(n2862), .B1(\REGISTERS[23][2] ), .B2(n2859), .ZN(n1578) );
  OAI221_X1 U1508 ( .B1(n2820), .B2(n1592), .C1(n2817), .C2(n1593), .A(n1594), 
        .ZN(n1583) );
  AOI22_X1 U1509 ( .A1(\REGISTERS[6][2] ), .A2(n2814), .B1(\REGISTERS[7][2] ), 
        .B2(n2811), .ZN(n1594) );
  OAI221_X1 U1510 ( .B1(n2868), .B2(n1542), .C1(n2865), .C2(n1543), .A(n1544), 
        .ZN(n1533) );
  AOI22_X1 U1511 ( .A1(\REGISTERS[22][3] ), .A2(n2862), .B1(\REGISTERS[23][3] ), .B2(n2859), .ZN(n1544) );
  OAI221_X1 U1512 ( .B1(n2820), .B2(n1558), .C1(n2817), .C2(n1559), .A(n1560), 
        .ZN(n1549) );
  AOI22_X1 U1513 ( .A1(\REGISTERS[6][3] ), .A2(n2814), .B1(\REGISTERS[7][3] ), 
        .B2(n2811), .ZN(n1560) );
  OAI221_X1 U1514 ( .B1(n2868), .B2(n1508), .C1(n2865), .C2(n1509), .A(n1510), 
        .ZN(n1499) );
  AOI22_X1 U1515 ( .A1(\REGISTERS[22][4] ), .A2(n2862), .B1(\REGISTERS[23][4] ), .B2(n2859), .ZN(n1510) );
  OAI221_X1 U1516 ( .B1(n2820), .B2(n1524), .C1(n2817), .C2(n1525), .A(n1526), 
        .ZN(n1515) );
  AOI22_X1 U1517 ( .A1(\REGISTERS[6][4] ), .A2(n2814), .B1(\REGISTERS[7][4] ), 
        .B2(n2811), .ZN(n1526) );
  OAI221_X1 U1518 ( .B1(n2868), .B2(n1474), .C1(n2865), .C2(n1475), .A(n1476), 
        .ZN(n1465) );
  AOI22_X1 U1519 ( .A1(\REGISTERS[22][5] ), .A2(n2862), .B1(\REGISTERS[23][5] ), .B2(n2859), .ZN(n1476) );
  OAI221_X1 U1520 ( .B1(n2820), .B2(n1490), .C1(n2817), .C2(n1491), .A(n1492), 
        .ZN(n1481) );
  AOI22_X1 U1521 ( .A1(\REGISTERS[6][5] ), .A2(n2814), .B1(\REGISTERS[7][5] ), 
        .B2(n2811), .ZN(n1492) );
  OAI221_X1 U1522 ( .B1(n2868), .B2(n1440), .C1(n2865), .C2(n1441), .A(n1442), 
        .ZN(n1431) );
  AOI22_X1 U1523 ( .A1(\REGISTERS[22][6] ), .A2(n2862), .B1(\REGISTERS[23][6] ), .B2(n2859), .ZN(n1442) );
  OAI221_X1 U1524 ( .B1(n2820), .B2(n1456), .C1(n2817), .C2(n1457), .A(n1458), 
        .ZN(n1447) );
  AOI22_X1 U1525 ( .A1(\REGISTERS[6][6] ), .A2(n2814), .B1(\REGISTERS[7][6] ), 
        .B2(n2811), .ZN(n1458) );
  OAI221_X1 U1526 ( .B1(n2868), .B2(n1406), .C1(n2865), .C2(n1407), .A(n1408), 
        .ZN(n1397) );
  AOI22_X1 U1527 ( .A1(\REGISTERS[22][7] ), .A2(n2862), .B1(\REGISTERS[23][7] ), .B2(n2859), .ZN(n1408) );
  OAI221_X1 U1528 ( .B1(n2820), .B2(n1422), .C1(n2817), .C2(n1423), .A(n1424), 
        .ZN(n1413) );
  AOI22_X1 U1529 ( .A1(\REGISTERS[6][7] ), .A2(n2814), .B1(\REGISTERS[7][7] ), 
        .B2(n2811), .ZN(n1424) );
  OAI221_X1 U1530 ( .B1(n2868), .B2(n1372), .C1(n2865), .C2(n1373), .A(n1374), 
        .ZN(n1363) );
  AOI22_X1 U1531 ( .A1(\REGISTERS[22][8] ), .A2(n2862), .B1(\REGISTERS[23][8] ), .B2(n2859), .ZN(n1374) );
  OAI221_X1 U1532 ( .B1(n2820), .B2(n1388), .C1(n2817), .C2(n1389), .A(n1390), 
        .ZN(n1379) );
  AOI22_X1 U1533 ( .A1(\REGISTERS[6][8] ), .A2(n2814), .B1(\REGISTERS[7][8] ), 
        .B2(n2811), .ZN(n1390) );
  OAI221_X1 U1534 ( .B1(n2868), .B2(n1338), .C1(n2865), .C2(n1339), .A(n1340), 
        .ZN(n1329) );
  AOI22_X1 U1535 ( .A1(\REGISTERS[22][9] ), .A2(n2862), .B1(\REGISTERS[23][9] ), .B2(n2859), .ZN(n1340) );
  OAI221_X1 U1536 ( .B1(n2820), .B2(n1354), .C1(n2817), .C2(n1355), .A(n1356), 
        .ZN(n1345) );
  AOI22_X1 U1537 ( .A1(\REGISTERS[6][9] ), .A2(n2814), .B1(\REGISTERS[7][9] ), 
        .B2(n2811), .ZN(n1356) );
  OAI221_X1 U1538 ( .B1(n2868), .B2(n1304), .C1(n2865), .C2(n1305), .A(n1306), 
        .ZN(n1295) );
  AOI22_X1 U1539 ( .A1(\REGISTERS[22][10] ), .A2(n2862), .B1(
        \REGISTERS[23][10] ), .B2(n2859), .ZN(n1306) );
  OAI221_X1 U1540 ( .B1(n2820), .B2(n1320), .C1(n2817), .C2(n1321), .A(n1322), 
        .ZN(n1311) );
  AOI22_X1 U1541 ( .A1(\REGISTERS[6][10] ), .A2(n2814), .B1(\REGISTERS[7][10] ), .B2(n2811), .ZN(n1322) );
  OAI221_X1 U1542 ( .B1(n2868), .B2(n1270), .C1(n2865), .C2(n1271), .A(n1272), 
        .ZN(n1261) );
  AOI22_X1 U1543 ( .A1(\REGISTERS[22][11] ), .A2(n2862), .B1(
        \REGISTERS[23][11] ), .B2(n2859), .ZN(n1272) );
  OAI221_X1 U1544 ( .B1(n2820), .B2(n1286), .C1(n2817), .C2(n1287), .A(n1288), 
        .ZN(n1277) );
  AOI22_X1 U1545 ( .A1(\REGISTERS[6][11] ), .A2(n2814), .B1(\REGISTERS[7][11] ), .B2(n2811), .ZN(n1288) );
  OAI221_X1 U1546 ( .B1(n2869), .B2(n1236), .C1(n2866), .C2(n1237), .A(n1238), 
        .ZN(n1227) );
  AOI22_X1 U1547 ( .A1(\REGISTERS[22][12] ), .A2(n2863), .B1(
        \REGISTERS[23][12] ), .B2(n2860), .ZN(n1238) );
  OAI221_X1 U1548 ( .B1(n2821), .B2(n1252), .C1(n2818), .C2(n1253), .A(n1254), 
        .ZN(n1243) );
  AOI22_X1 U1549 ( .A1(\REGISTERS[6][12] ), .A2(n2815), .B1(\REGISTERS[7][12] ), .B2(n2812), .ZN(n1254) );
  OAI221_X1 U1550 ( .B1(n2869), .B2(n1202), .C1(n2866), .C2(n1203), .A(n1204), 
        .ZN(n1193) );
  AOI22_X1 U1551 ( .A1(\REGISTERS[22][13] ), .A2(n2863), .B1(
        \REGISTERS[23][13] ), .B2(n2860), .ZN(n1204) );
  OAI221_X1 U1552 ( .B1(n2821), .B2(n1218), .C1(n2818), .C2(n1219), .A(n1220), 
        .ZN(n1209) );
  AOI22_X1 U1553 ( .A1(\REGISTERS[6][13] ), .A2(n2815), .B1(\REGISTERS[7][13] ), .B2(n2812), .ZN(n1220) );
  OAI221_X1 U1554 ( .B1(n2869), .B2(n1168), .C1(n2866), .C2(n1169), .A(n1170), 
        .ZN(n1159) );
  AOI22_X1 U1555 ( .A1(\REGISTERS[22][14] ), .A2(n2863), .B1(
        \REGISTERS[23][14] ), .B2(n2860), .ZN(n1170) );
  OAI221_X1 U1556 ( .B1(n2821), .B2(n1184), .C1(n2818), .C2(n1185), .A(n1186), 
        .ZN(n1175) );
  AOI22_X1 U1557 ( .A1(\REGISTERS[6][14] ), .A2(n2815), .B1(\REGISTERS[7][14] ), .B2(n2812), .ZN(n1186) );
  OAI221_X1 U1558 ( .B1(n2869), .B2(n1134), .C1(n2866), .C2(n1135), .A(n1136), 
        .ZN(n1125) );
  AOI22_X1 U1559 ( .A1(\REGISTERS[22][15] ), .A2(n2863), .B1(
        \REGISTERS[23][15] ), .B2(n2860), .ZN(n1136) );
  OAI221_X1 U1560 ( .B1(n2821), .B2(n1150), .C1(n2818), .C2(n1151), .A(n1152), 
        .ZN(n1141) );
  AOI22_X1 U1561 ( .A1(\REGISTERS[6][15] ), .A2(n2815), .B1(\REGISTERS[7][15] ), .B2(n2812), .ZN(n1152) );
  OAI221_X1 U1562 ( .B1(n2869), .B2(n1100), .C1(n2866), .C2(n1101), .A(n1102), 
        .ZN(n1091) );
  AOI22_X1 U1563 ( .A1(\REGISTERS[22][16] ), .A2(n2863), .B1(
        \REGISTERS[23][16] ), .B2(n2860), .ZN(n1102) );
  OAI221_X1 U1564 ( .B1(n2821), .B2(n1116), .C1(n2818), .C2(n1117), .A(n1118), 
        .ZN(n1107) );
  AOI22_X1 U1565 ( .A1(\REGISTERS[6][16] ), .A2(n2815), .B1(\REGISTERS[7][16] ), .B2(n2812), .ZN(n1118) );
  OAI221_X1 U1566 ( .B1(n2869), .B2(n1066), .C1(n2866), .C2(n1067), .A(n1068), 
        .ZN(n1057) );
  AOI22_X1 U1567 ( .A1(\REGISTERS[22][17] ), .A2(n2863), .B1(
        \REGISTERS[23][17] ), .B2(n2860), .ZN(n1068) );
  OAI221_X1 U1568 ( .B1(n2821), .B2(n1082), .C1(n2818), .C2(n1083), .A(n1084), 
        .ZN(n1073) );
  AOI22_X1 U1569 ( .A1(\REGISTERS[6][17] ), .A2(n2815), .B1(\REGISTERS[7][17] ), .B2(n2812), .ZN(n1084) );
  OAI221_X1 U1570 ( .B1(n2869), .B2(n1032), .C1(n2866), .C2(n1033), .A(n1034), 
        .ZN(n1023) );
  AOI22_X1 U1571 ( .A1(\REGISTERS[22][18] ), .A2(n2863), .B1(
        \REGISTERS[23][18] ), .B2(n2860), .ZN(n1034) );
  OAI221_X1 U1572 ( .B1(n2821), .B2(n1048), .C1(n2818), .C2(n1049), .A(n1050), 
        .ZN(n1039) );
  AOI22_X1 U1573 ( .A1(\REGISTERS[6][18] ), .A2(n2815), .B1(\REGISTERS[7][18] ), .B2(n2812), .ZN(n1050) );
  OAI221_X1 U1574 ( .B1(n2869), .B2(n998), .C1(n2866), .C2(n999), .A(n1000), 
        .ZN(n989) );
  AOI22_X1 U1575 ( .A1(\REGISTERS[22][19] ), .A2(n2863), .B1(
        \REGISTERS[23][19] ), .B2(n2860), .ZN(n1000) );
  OAI221_X1 U1576 ( .B1(n2821), .B2(n1014), .C1(n2818), .C2(n1015), .A(n1016), 
        .ZN(n1005) );
  AOI22_X1 U1577 ( .A1(\REGISTERS[6][19] ), .A2(n2815), .B1(\REGISTERS[7][19] ), .B2(n2812), .ZN(n1016) );
  OAI221_X1 U1578 ( .B1(n2869), .B2(n964), .C1(n2866), .C2(n965), .A(n966), 
        .ZN(n955) );
  AOI22_X1 U1579 ( .A1(\REGISTERS[22][20] ), .A2(n2863), .B1(
        \REGISTERS[23][20] ), .B2(n2860), .ZN(n966) );
  OAI221_X1 U1580 ( .B1(n2821), .B2(n980), .C1(n2818), .C2(n981), .A(n982), 
        .ZN(n971) );
  AOI22_X1 U1581 ( .A1(\REGISTERS[6][20] ), .A2(n2815), .B1(\REGISTERS[7][20] ), .B2(n2812), .ZN(n982) );
  OAI221_X1 U1582 ( .B1(n2869), .B2(n930), .C1(n2866), .C2(n931), .A(n932), 
        .ZN(n921) );
  AOI22_X1 U1583 ( .A1(\REGISTERS[22][21] ), .A2(n2863), .B1(
        \REGISTERS[23][21] ), .B2(n2860), .ZN(n932) );
  OAI221_X1 U1584 ( .B1(n2821), .B2(n946), .C1(n2818), .C2(n947), .A(n948), 
        .ZN(n937) );
  AOI22_X1 U1585 ( .A1(\REGISTERS[6][21] ), .A2(n2815), .B1(\REGISTERS[7][21] ), .B2(n2812), .ZN(n948) );
  OAI221_X1 U1586 ( .B1(n2869), .B2(n896), .C1(n2866), .C2(n897), .A(n898), 
        .ZN(n887) );
  AOI22_X1 U1587 ( .A1(\REGISTERS[22][22] ), .A2(n2863), .B1(
        \REGISTERS[23][22] ), .B2(n2860), .ZN(n898) );
  OAI221_X1 U1588 ( .B1(n2821), .B2(n912), .C1(n2818), .C2(n913), .A(n914), 
        .ZN(n903) );
  AOI22_X1 U1589 ( .A1(\REGISTERS[6][22] ), .A2(n2815), .B1(\REGISTERS[7][22] ), .B2(n2812), .ZN(n914) );
  OAI221_X1 U1590 ( .B1(n2869), .B2(n862), .C1(n2866), .C2(n863), .A(n864), 
        .ZN(n853) );
  AOI22_X1 U1591 ( .A1(\REGISTERS[22][23] ), .A2(n2863), .B1(
        \REGISTERS[23][23] ), .B2(n2860), .ZN(n864) );
  OAI221_X1 U1592 ( .B1(n2821), .B2(n878), .C1(n2818), .C2(n879), .A(n880), 
        .ZN(n869) );
  AOI22_X1 U1593 ( .A1(\REGISTERS[6][23] ), .A2(n2815), .B1(\REGISTERS[7][23] ), .B2(n2812), .ZN(n880) );
  OAI221_X1 U1594 ( .B1(n1656), .B2(n2760), .C1(n1657), .C2(n2757), .A(n2290), 
        .ZN(n2274) );
  AOI22_X1 U1595 ( .A1(n2754), .A2(\REGISTERS[18][0] ), .B1(n2753), .B2(
        \REGISTERS[19][0] ), .ZN(n2290) );
  OAI221_X1 U1596 ( .B1(n1613), .B2(n2760), .C1(n1614), .C2(n2757), .A(n2263), 
        .ZN(n2256) );
  AOI22_X1 U1597 ( .A1(n2754), .A2(\REGISTERS[18][1] ), .B1(n2753), .B2(
        \REGISTERS[19][1] ), .ZN(n2263) );
  OAI221_X1 U1598 ( .B1(n1579), .B2(n2760), .C1(n1580), .C2(n2757), .A(n2245), 
        .ZN(n2238) );
  AOI22_X1 U1599 ( .A1(n2754), .A2(\REGISTERS[18][2] ), .B1(n2753), .B2(
        \REGISTERS[19][2] ), .ZN(n2245) );
  OAI221_X1 U1600 ( .B1(n1545), .B2(n2760), .C1(n1546), .C2(n2757), .A(n2227), 
        .ZN(n2220) );
  AOI22_X1 U1601 ( .A1(n2754), .A2(\REGISTERS[18][3] ), .B1(n2753), .B2(
        \REGISTERS[19][3] ), .ZN(n2227) );
  OAI221_X1 U1602 ( .B1(n1511), .B2(n2760), .C1(n1512), .C2(n2757), .A(n2209), 
        .ZN(n2202) );
  AOI22_X1 U1603 ( .A1(n2754), .A2(\REGISTERS[18][4] ), .B1(n2753), .B2(
        \REGISTERS[19][4] ), .ZN(n2209) );
  OAI221_X1 U1604 ( .B1(n1477), .B2(n2760), .C1(n1478), .C2(n2757), .A(n2191), 
        .ZN(n2184) );
  AOI22_X1 U1605 ( .A1(n2754), .A2(\REGISTERS[18][5] ), .B1(n2753), .B2(
        \REGISTERS[19][5] ), .ZN(n2191) );
  OAI221_X1 U1606 ( .B1(n1443), .B2(n2760), .C1(n1444), .C2(n2757), .A(n2173), 
        .ZN(n2166) );
  AOI22_X1 U1607 ( .A1(n2754), .A2(\REGISTERS[18][6] ), .B1(n2753), .B2(
        \REGISTERS[19][6] ), .ZN(n2173) );
  OAI221_X1 U1608 ( .B1(n1409), .B2(n2760), .C1(n1410), .C2(n2757), .A(n2155), 
        .ZN(n2148) );
  AOI22_X1 U1609 ( .A1(n2754), .A2(\REGISTERS[18][7] ), .B1(n2753), .B2(
        \REGISTERS[19][7] ), .ZN(n2155) );
  OAI221_X1 U1610 ( .B1(n1375), .B2(n2760), .C1(n1376), .C2(n2757), .A(n2137), 
        .ZN(n2130) );
  AOI22_X1 U1611 ( .A1(n2754), .A2(\REGISTERS[18][8] ), .B1(n2752), .B2(
        \REGISTERS[19][8] ), .ZN(n2137) );
  OAI221_X1 U1612 ( .B1(n1341), .B2(n2760), .C1(n1342), .C2(n2757), .A(n2119), 
        .ZN(n2112) );
  AOI22_X1 U1613 ( .A1(n2754), .A2(\REGISTERS[18][9] ), .B1(n2752), .B2(
        \REGISTERS[19][9] ), .ZN(n2119) );
  OAI221_X1 U1614 ( .B1(n1307), .B2(n2760), .C1(n1308), .C2(n2757), .A(n2101), 
        .ZN(n2094) );
  AOI22_X1 U1615 ( .A1(n2754), .A2(\REGISTERS[18][10] ), .B1(n2752), .B2(
        \REGISTERS[19][10] ), .ZN(n2101) );
  OAI221_X1 U1616 ( .B1(n1273), .B2(n2760), .C1(n1274), .C2(n2757), .A(n2083), 
        .ZN(n2076) );
  AOI22_X1 U1617 ( .A1(n2754), .A2(\REGISTERS[18][11] ), .B1(n2752), .B2(
        \REGISTERS[19][11] ), .ZN(n2083) );
  OAI221_X1 U1618 ( .B1(n1239), .B2(n2761), .C1(n1240), .C2(n2758), .A(n2065), 
        .ZN(n2058) );
  AOI22_X1 U1619 ( .A1(n2755), .A2(\REGISTERS[18][12] ), .B1(n2752), .B2(
        \REGISTERS[19][12] ), .ZN(n2065) );
  OAI221_X1 U1620 ( .B1(n1205), .B2(n2761), .C1(n1206), .C2(n2758), .A(n2047), 
        .ZN(n2040) );
  AOI22_X1 U1621 ( .A1(n2755), .A2(\REGISTERS[18][13] ), .B1(n2752), .B2(
        \REGISTERS[19][13] ), .ZN(n2047) );
  OAI221_X1 U1622 ( .B1(n1171), .B2(n2761), .C1(n1172), .C2(n2758), .A(n2029), 
        .ZN(n2022) );
  AOI22_X1 U1623 ( .A1(n2755), .A2(\REGISTERS[18][14] ), .B1(n2752), .B2(
        \REGISTERS[19][14] ), .ZN(n2029) );
  OAI221_X1 U1624 ( .B1(n1137), .B2(n2761), .C1(n1138), .C2(n2758), .A(n2011), 
        .ZN(n2004) );
  AOI22_X1 U1625 ( .A1(n2755), .A2(\REGISTERS[18][15] ), .B1(n2752), .B2(
        \REGISTERS[19][15] ), .ZN(n2011) );
  OAI221_X1 U1626 ( .B1(n1103), .B2(n2761), .C1(n1104), .C2(n2758), .A(n1993), 
        .ZN(n1986) );
  AOI22_X1 U1627 ( .A1(n2755), .A2(\REGISTERS[18][16] ), .B1(n2752), .B2(
        \REGISTERS[19][16] ), .ZN(n1993) );
  OAI221_X1 U1628 ( .B1(n1069), .B2(n2761), .C1(n1070), .C2(n2758), .A(n1975), 
        .ZN(n1968) );
  AOI22_X1 U1629 ( .A1(n2755), .A2(\REGISTERS[18][17] ), .B1(n2752), .B2(
        \REGISTERS[19][17] ), .ZN(n1975) );
  OAI221_X1 U1630 ( .B1(n1035), .B2(n2761), .C1(n1036), .C2(n2758), .A(n1957), 
        .ZN(n1950) );
  AOI22_X1 U1631 ( .A1(n2755), .A2(\REGISTERS[18][18] ), .B1(n2752), .B2(
        \REGISTERS[19][18] ), .ZN(n1957) );
  OAI221_X1 U1632 ( .B1(n1001), .B2(n2761), .C1(n1002), .C2(n2758), .A(n1939), 
        .ZN(n1932) );
  AOI22_X1 U1633 ( .A1(n2755), .A2(\REGISTERS[18][19] ), .B1(n2752), .B2(
        \REGISTERS[19][19] ), .ZN(n1939) );
  OAI221_X1 U1634 ( .B1(n967), .B2(n2761), .C1(n968), .C2(n2758), .A(n1921), 
        .ZN(n1914) );
  AOI22_X1 U1635 ( .A1(n2755), .A2(\REGISTERS[18][20] ), .B1(n2751), .B2(
        \REGISTERS[19][20] ), .ZN(n1921) );
  OAI221_X1 U1636 ( .B1(n933), .B2(n2761), .C1(n934), .C2(n2758), .A(n1903), 
        .ZN(n1896) );
  AOI22_X1 U1637 ( .A1(n2755), .A2(\REGISTERS[18][21] ), .B1(n2751), .B2(
        \REGISTERS[19][21] ), .ZN(n1903) );
  OAI221_X1 U1638 ( .B1(n899), .B2(n2761), .C1(n900), .C2(n2758), .A(n1885), 
        .ZN(n1878) );
  AOI22_X1 U1639 ( .A1(n2755), .A2(\REGISTERS[18][22] ), .B1(n2751), .B2(
        \REGISTERS[19][22] ), .ZN(n1885) );
  OAI221_X1 U1640 ( .B1(n865), .B2(n2761), .C1(n866), .C2(n2758), .A(n1867), 
        .ZN(n1860) );
  AOI22_X1 U1641 ( .A1(n2755), .A2(\REGISTERS[18][23] ), .B1(n2751), .B2(
        \REGISTERS[19][23] ), .ZN(n1867) );
  OAI221_X1 U1642 ( .B1(n2856), .B2(n1656), .C1(n2853), .C2(n1657), .A(n1658), 
        .ZN(n1634) );
  AOI22_X1 U1643 ( .A1(\REGISTERS[18][0] ), .A2(n2850), .B1(\REGISTERS[19][0] ), .B2(n2847), .ZN(n1658) );
  OAI221_X1 U1644 ( .B1(n2856), .B2(n1613), .C1(n2853), .C2(n1614), .A(n1615), 
        .ZN(n1600) );
  AOI22_X1 U1645 ( .A1(\REGISTERS[18][1] ), .A2(n2850), .B1(\REGISTERS[19][1] ), .B2(n2847), .ZN(n1615) );
  OAI221_X1 U1646 ( .B1(n2856), .B2(n1579), .C1(n2853), .C2(n1580), .A(n1581), 
        .ZN(n1566) );
  AOI22_X1 U1647 ( .A1(\REGISTERS[18][2] ), .A2(n2850), .B1(\REGISTERS[19][2] ), .B2(n2847), .ZN(n1581) );
  OAI221_X1 U1648 ( .B1(n2856), .B2(n1545), .C1(n2853), .C2(n1546), .A(n1547), 
        .ZN(n1532) );
  AOI22_X1 U1649 ( .A1(\REGISTERS[18][3] ), .A2(n2850), .B1(\REGISTERS[19][3] ), .B2(n2847), .ZN(n1547) );
  OAI221_X1 U1650 ( .B1(n2856), .B2(n1511), .C1(n2853), .C2(n1512), .A(n1513), 
        .ZN(n1498) );
  AOI22_X1 U1651 ( .A1(\REGISTERS[18][4] ), .A2(n2850), .B1(\REGISTERS[19][4] ), .B2(n2847), .ZN(n1513) );
  OAI221_X1 U1652 ( .B1(n2856), .B2(n1477), .C1(n2853), .C2(n1478), .A(n1479), 
        .ZN(n1464) );
  AOI22_X1 U1653 ( .A1(\REGISTERS[18][5] ), .A2(n2850), .B1(\REGISTERS[19][5] ), .B2(n2847), .ZN(n1479) );
  OAI221_X1 U1654 ( .B1(n2856), .B2(n1443), .C1(n2853), .C2(n1444), .A(n1445), 
        .ZN(n1430) );
  AOI22_X1 U1655 ( .A1(\REGISTERS[18][6] ), .A2(n2850), .B1(\REGISTERS[19][6] ), .B2(n2847), .ZN(n1445) );
  OAI221_X1 U1656 ( .B1(n2856), .B2(n1409), .C1(n2853), .C2(n1410), .A(n1411), 
        .ZN(n1396) );
  AOI22_X1 U1657 ( .A1(\REGISTERS[18][7] ), .A2(n2850), .B1(\REGISTERS[19][7] ), .B2(n2847), .ZN(n1411) );
  OAI221_X1 U1658 ( .B1(n2856), .B2(n1375), .C1(n2853), .C2(n1376), .A(n1377), 
        .ZN(n1362) );
  AOI22_X1 U1659 ( .A1(\REGISTERS[18][8] ), .A2(n2850), .B1(\REGISTERS[19][8] ), .B2(n2847), .ZN(n1377) );
  OAI221_X1 U1660 ( .B1(n2856), .B2(n1341), .C1(n2853), .C2(n1342), .A(n1343), 
        .ZN(n1328) );
  AOI22_X1 U1661 ( .A1(\REGISTERS[18][9] ), .A2(n2850), .B1(\REGISTERS[19][9] ), .B2(n2847), .ZN(n1343) );
  OAI221_X1 U1662 ( .B1(n2856), .B2(n1307), .C1(n2853), .C2(n1308), .A(n1309), 
        .ZN(n1294) );
  AOI22_X1 U1663 ( .A1(\REGISTERS[18][10] ), .A2(n2850), .B1(
        \REGISTERS[19][10] ), .B2(n2847), .ZN(n1309) );
  OAI221_X1 U1664 ( .B1(n2856), .B2(n1273), .C1(n2853), .C2(n1274), .A(n1275), 
        .ZN(n1260) );
  AOI22_X1 U1665 ( .A1(\REGISTERS[18][11] ), .A2(n2850), .B1(
        \REGISTERS[19][11] ), .B2(n2847), .ZN(n1275) );
  OAI221_X1 U1666 ( .B1(n2857), .B2(n1239), .C1(n2854), .C2(n1240), .A(n1241), 
        .ZN(n1226) );
  AOI22_X1 U1667 ( .A1(\REGISTERS[18][12] ), .A2(n2851), .B1(
        \REGISTERS[19][12] ), .B2(n2848), .ZN(n1241) );
  OAI221_X1 U1668 ( .B1(n2857), .B2(n1205), .C1(n2854), .C2(n1206), .A(n1207), 
        .ZN(n1192) );
  AOI22_X1 U1669 ( .A1(\REGISTERS[18][13] ), .A2(n2851), .B1(
        \REGISTERS[19][13] ), .B2(n2848), .ZN(n1207) );
  OAI221_X1 U1670 ( .B1(n2857), .B2(n1171), .C1(n2854), .C2(n1172), .A(n1173), 
        .ZN(n1158) );
  AOI22_X1 U1671 ( .A1(\REGISTERS[18][14] ), .A2(n2851), .B1(
        \REGISTERS[19][14] ), .B2(n2848), .ZN(n1173) );
  OAI221_X1 U1672 ( .B1(n2857), .B2(n1137), .C1(n2854), .C2(n1138), .A(n1139), 
        .ZN(n1124) );
  AOI22_X1 U1673 ( .A1(\REGISTERS[18][15] ), .A2(n2851), .B1(
        \REGISTERS[19][15] ), .B2(n2848), .ZN(n1139) );
  OAI221_X1 U1674 ( .B1(n2857), .B2(n1103), .C1(n2854), .C2(n1104), .A(n1105), 
        .ZN(n1090) );
  AOI22_X1 U1675 ( .A1(\REGISTERS[18][16] ), .A2(n2851), .B1(
        \REGISTERS[19][16] ), .B2(n2848), .ZN(n1105) );
  OAI221_X1 U1676 ( .B1(n2857), .B2(n1069), .C1(n2854), .C2(n1070), .A(n1071), 
        .ZN(n1056) );
  AOI22_X1 U1677 ( .A1(\REGISTERS[18][17] ), .A2(n2851), .B1(
        \REGISTERS[19][17] ), .B2(n2848), .ZN(n1071) );
  OAI221_X1 U1678 ( .B1(n2857), .B2(n1035), .C1(n2854), .C2(n1036), .A(n1037), 
        .ZN(n1022) );
  AOI22_X1 U1679 ( .A1(\REGISTERS[18][18] ), .A2(n2851), .B1(
        \REGISTERS[19][18] ), .B2(n2848), .ZN(n1037) );
  OAI221_X1 U1680 ( .B1(n2857), .B2(n1001), .C1(n2854), .C2(n1002), .A(n1003), 
        .ZN(n988) );
  AOI22_X1 U1681 ( .A1(\REGISTERS[18][19] ), .A2(n2851), .B1(
        \REGISTERS[19][19] ), .B2(n2848), .ZN(n1003) );
  OAI221_X1 U1682 ( .B1(n2857), .B2(n967), .C1(n2854), .C2(n968), .A(n969), 
        .ZN(n954) );
  AOI22_X1 U1683 ( .A1(\REGISTERS[18][20] ), .A2(n2851), .B1(
        \REGISTERS[19][20] ), .B2(n2848), .ZN(n969) );
  OAI221_X1 U1684 ( .B1(n2857), .B2(n933), .C1(n2854), .C2(n934), .A(n935), 
        .ZN(n920) );
  AOI22_X1 U1685 ( .A1(\REGISTERS[18][21] ), .A2(n2851), .B1(
        \REGISTERS[19][21] ), .B2(n2848), .ZN(n935) );
  OAI221_X1 U1686 ( .B1(n2857), .B2(n899), .C1(n2854), .C2(n900), .A(n901), 
        .ZN(n886) );
  AOI22_X1 U1687 ( .A1(\REGISTERS[18][22] ), .A2(n2851), .B1(
        \REGISTERS[19][22] ), .B2(n2848), .ZN(n901) );
  OAI221_X1 U1688 ( .B1(n2857), .B2(n865), .C1(n2854), .C2(n866), .A(n867), 
        .ZN(n852) );
  AOI22_X1 U1689 ( .A1(\REGISTERS[18][23] ), .A2(n2851), .B1(
        \REGISTERS[19][23] ), .B2(n2848), .ZN(n867) );
  AOI22_X1 U1690 ( .A1(\REGISTERS[2][24] ), .A2(n2804), .B1(\REGISTERS[3][24] ), .B2(n2801), .ZN(n849) );
  AOI22_X1 U1691 ( .A1(\REGISTERS[2][25] ), .A2(n2804), .B1(\REGISTERS[3][25] ), .B2(n2801), .ZN(n815) );
  AOI22_X1 U1692 ( .A1(\REGISTERS[2][26] ), .A2(n2804), .B1(\REGISTERS[3][26] ), .B2(n2801), .ZN(n781) );
  AOI22_X1 U1693 ( .A1(\REGISTERS[2][27] ), .A2(n2804), .B1(\REGISTERS[3][27] ), .B2(n2801), .ZN(n747) );
  AOI22_X1 U1694 ( .A1(\REGISTERS[2][28] ), .A2(n2804), .B1(\REGISTERS[3][28] ), .B2(n2801), .ZN(n713) );
  AOI22_X1 U1695 ( .A1(\REGISTERS[2][29] ), .A2(n2804), .B1(\REGISTERS[3][29] ), .B2(n2801), .ZN(n679) );
  AOI22_X1 U1696 ( .A1(\REGISTERS[2][30] ), .A2(n2804), .B1(\REGISTERS[3][30] ), .B2(n2801), .ZN(n645) );
  AOI22_X1 U1697 ( .A1(\REGISTERS[2][31] ), .A2(n2804), .B1(\REGISTERS[3][31] ), .B2(n2801), .ZN(n609) );
  AOI22_X1 U1698 ( .A1(n2706), .A2(\REGISTERS[2][0] ), .B1(n2705), .B2(
        \REGISTERS[3][0] ), .ZN(n2304) );
  AOI22_X1 U1699 ( .A1(n2706), .A2(\REGISTERS[2][1] ), .B1(n2705), .B2(
        \REGISTERS[3][1] ), .ZN(n2271) );
  AOI22_X1 U1700 ( .A1(n2706), .A2(\REGISTERS[2][2] ), .B1(n2705), .B2(
        \REGISTERS[3][2] ), .ZN(n2253) );
  AOI22_X1 U1701 ( .A1(n2706), .A2(\REGISTERS[2][3] ), .B1(n2705), .B2(
        \REGISTERS[3][3] ), .ZN(n2235) );
  AOI22_X1 U1702 ( .A1(n2706), .A2(\REGISTERS[2][4] ), .B1(n2705), .B2(
        \REGISTERS[3][4] ), .ZN(n2217) );
  AOI22_X1 U1703 ( .A1(n2706), .A2(\REGISTERS[2][5] ), .B1(n2705), .B2(
        \REGISTERS[3][5] ), .ZN(n2199) );
  AOI22_X1 U1704 ( .A1(n2706), .A2(\REGISTERS[2][6] ), .B1(n2705), .B2(
        \REGISTERS[3][6] ), .ZN(n2181) );
  AOI22_X1 U1705 ( .A1(n2706), .A2(\REGISTERS[2][7] ), .B1(n2705), .B2(
        \REGISTERS[3][7] ), .ZN(n2163) );
  AOI22_X1 U1706 ( .A1(n2706), .A2(\REGISTERS[2][8] ), .B1(n2704), .B2(
        \REGISTERS[3][8] ), .ZN(n2145) );
  AOI22_X1 U1707 ( .A1(n2706), .A2(\REGISTERS[2][9] ), .B1(n2704), .B2(
        \REGISTERS[3][9] ), .ZN(n2127) );
  AOI22_X1 U1708 ( .A1(n2706), .A2(\REGISTERS[2][10] ), .B1(n2704), .B2(
        \REGISTERS[3][10] ), .ZN(n2109) );
  AOI22_X1 U1709 ( .A1(n2706), .A2(\REGISTERS[2][11] ), .B1(n2704), .B2(
        \REGISTERS[3][11] ), .ZN(n2091) );
  AOI22_X1 U1710 ( .A1(n2707), .A2(\REGISTERS[2][12] ), .B1(n2704), .B2(
        \REGISTERS[3][12] ), .ZN(n2073) );
  AOI22_X1 U1711 ( .A1(n2707), .A2(\REGISTERS[2][13] ), .B1(n2704), .B2(
        \REGISTERS[3][13] ), .ZN(n2055) );
  AOI22_X1 U1712 ( .A1(n2707), .A2(\REGISTERS[2][14] ), .B1(n2704), .B2(
        \REGISTERS[3][14] ), .ZN(n2037) );
  AOI22_X1 U1713 ( .A1(n2707), .A2(\REGISTERS[2][15] ), .B1(n2704), .B2(
        \REGISTERS[3][15] ), .ZN(n2019) );
  AOI22_X1 U1714 ( .A1(n2707), .A2(\REGISTERS[2][16] ), .B1(n2704), .B2(
        \REGISTERS[3][16] ), .ZN(n2001) );
  AOI22_X1 U1715 ( .A1(n2707), .A2(\REGISTERS[2][17] ), .B1(n2704), .B2(
        \REGISTERS[3][17] ), .ZN(n1983) );
  AOI22_X1 U1716 ( .A1(n2707), .A2(\REGISTERS[2][18] ), .B1(n2704), .B2(
        \REGISTERS[3][18] ), .ZN(n1965) );
  AOI22_X1 U1717 ( .A1(n2707), .A2(\REGISTERS[2][19] ), .B1(n2704), .B2(
        \REGISTERS[3][19] ), .ZN(n1947) );
  AOI22_X1 U1718 ( .A1(n2707), .A2(\REGISTERS[2][20] ), .B1(n2703), .B2(
        \REGISTERS[3][20] ), .ZN(n1929) );
  AOI22_X1 U1719 ( .A1(n2707), .A2(\REGISTERS[2][21] ), .B1(n2703), .B2(
        \REGISTERS[3][21] ), .ZN(n1911) );
  AOI22_X1 U1720 ( .A1(n2707), .A2(\REGISTERS[2][22] ), .B1(n2703), .B2(
        \REGISTERS[3][22] ), .ZN(n1893) );
  AOI22_X1 U1721 ( .A1(n2707), .A2(\REGISTERS[2][23] ), .B1(n2703), .B2(
        \REGISTERS[3][23] ), .ZN(n1875) );
  AOI22_X1 U1722 ( .A1(n2708), .A2(\REGISTERS[2][24] ), .B1(n2703), .B2(
        \REGISTERS[3][24] ), .ZN(n1857) );
  AOI22_X1 U1723 ( .A1(n2708), .A2(\REGISTERS[2][25] ), .B1(n2703), .B2(
        \REGISTERS[3][25] ), .ZN(n1839) );
  AOI22_X1 U1724 ( .A1(n2708), .A2(\REGISTERS[2][26] ), .B1(n2703), .B2(
        \REGISTERS[3][26] ), .ZN(n1821) );
  AOI22_X1 U1725 ( .A1(n2708), .A2(\REGISTERS[2][27] ), .B1(n2703), .B2(
        \REGISTERS[3][27] ), .ZN(n1803) );
  AOI22_X1 U1726 ( .A1(n2708), .A2(\REGISTERS[2][28] ), .B1(n2703), .B2(
        \REGISTERS[3][28] ), .ZN(n1785) );
  AOI22_X1 U1727 ( .A1(n2708), .A2(\REGISTERS[2][29] ), .B1(n2703), .B2(
        \REGISTERS[3][29] ), .ZN(n1767) );
  AOI22_X1 U1728 ( .A1(n2708), .A2(\REGISTERS[2][30] ), .B1(n2703), .B2(
        \REGISTERS[3][30] ), .ZN(n1749) );
  AOI22_X1 U1729 ( .A1(n2708), .A2(\REGISTERS[2][31] ), .B1(n2703), .B2(
        \REGISTERS[3][31] ), .ZN(n1729) );
  AOI22_X1 U1730 ( .A1(\REGISTERS[2][0] ), .A2(n2802), .B1(\REGISTERS[3][0] ), 
        .B2(n2799), .ZN(n1680) );
  AOI22_X1 U1731 ( .A1(\REGISTERS[2][1] ), .A2(n2802), .B1(\REGISTERS[3][1] ), 
        .B2(n2799), .ZN(n1631) );
  AOI22_X1 U1732 ( .A1(\REGISTERS[2][2] ), .A2(n2802), .B1(\REGISTERS[3][2] ), 
        .B2(n2799), .ZN(n1597) );
  AOI22_X1 U1733 ( .A1(\REGISTERS[2][3] ), .A2(n2802), .B1(\REGISTERS[3][3] ), 
        .B2(n2799), .ZN(n1563) );
  AOI22_X1 U1734 ( .A1(\REGISTERS[2][4] ), .A2(n2802), .B1(\REGISTERS[3][4] ), 
        .B2(n2799), .ZN(n1529) );
  AOI22_X1 U1735 ( .A1(\REGISTERS[2][5] ), .A2(n2802), .B1(\REGISTERS[3][5] ), 
        .B2(n2799), .ZN(n1495) );
  AOI22_X1 U1736 ( .A1(\REGISTERS[2][6] ), .A2(n2802), .B1(\REGISTERS[3][6] ), 
        .B2(n2799), .ZN(n1461) );
  AOI22_X1 U1737 ( .A1(\REGISTERS[2][7] ), .A2(n2802), .B1(\REGISTERS[3][7] ), 
        .B2(n2799), .ZN(n1427) );
  AOI22_X1 U1738 ( .A1(\REGISTERS[2][8] ), .A2(n2802), .B1(\REGISTERS[3][8] ), 
        .B2(n2799), .ZN(n1393) );
  AOI22_X1 U1739 ( .A1(\REGISTERS[2][9] ), .A2(n2802), .B1(\REGISTERS[3][9] ), 
        .B2(n2799), .ZN(n1359) );
  AOI22_X1 U1740 ( .A1(\REGISTERS[2][10] ), .A2(n2802), .B1(\REGISTERS[3][10] ), .B2(n2799), .ZN(n1325) );
  AOI22_X1 U1741 ( .A1(\REGISTERS[2][11] ), .A2(n2802), .B1(\REGISTERS[3][11] ), .B2(n2799), .ZN(n1291) );
  AOI22_X1 U1742 ( .A1(\REGISTERS[2][12] ), .A2(n2803), .B1(\REGISTERS[3][12] ), .B2(n2800), .ZN(n1257) );
  AOI22_X1 U1743 ( .A1(\REGISTERS[2][13] ), .A2(n2803), .B1(\REGISTERS[3][13] ), .B2(n2800), .ZN(n1223) );
  AOI22_X1 U1744 ( .A1(\REGISTERS[2][14] ), .A2(n2803), .B1(\REGISTERS[3][14] ), .B2(n2800), .ZN(n1189) );
  AOI22_X1 U1745 ( .A1(\REGISTERS[2][15] ), .A2(n2803), .B1(\REGISTERS[3][15] ), .B2(n2800), .ZN(n1155) );
  AOI22_X1 U1746 ( .A1(\REGISTERS[2][16] ), .A2(n2803), .B1(\REGISTERS[3][16] ), .B2(n2800), .ZN(n1121) );
  AOI22_X1 U1747 ( .A1(\REGISTERS[2][17] ), .A2(n2803), .B1(\REGISTERS[3][17] ), .B2(n2800), .ZN(n1087) );
  AOI22_X1 U1748 ( .A1(\REGISTERS[2][18] ), .A2(n2803), .B1(\REGISTERS[3][18] ), .B2(n2800), .ZN(n1053) );
  AOI22_X1 U1749 ( .A1(\REGISTERS[2][19] ), .A2(n2803), .B1(\REGISTERS[3][19] ), .B2(n2800), .ZN(n1019) );
  AOI22_X1 U1750 ( .A1(\REGISTERS[2][20] ), .A2(n2803), .B1(\REGISTERS[3][20] ), .B2(n2800), .ZN(n985) );
  AOI22_X1 U1751 ( .A1(\REGISTERS[2][21] ), .A2(n2803), .B1(\REGISTERS[3][21] ), .B2(n2800), .ZN(n951) );
  AOI22_X1 U1752 ( .A1(\REGISTERS[2][22] ), .A2(n2803), .B1(\REGISTERS[3][22] ), .B2(n2800), .ZN(n917) );
  AOI22_X1 U1753 ( .A1(\REGISTERS[2][23] ), .A2(n2803), .B1(\REGISTERS[3][23] ), .B2(n2800), .ZN(n883) );
  AND3_X1 U1754 ( .A1(n3099), .A2(n2305), .A3(ADD_RD1[1]), .ZN(n2284) );
  AND3_X1 U1755 ( .A1(n3099), .A2(n1681), .A3(ADD_RD2[1]), .ZN(n1648) );
  AND3_X1 U1756 ( .A1(ADD_RD2[1]), .A2(n3099), .A3(ADD_RD2[2]), .ZN(n1642) );
  AND3_X1 U1757 ( .A1(ADD_RD1[1]), .A2(n3099), .A3(ADD_RD1[2]), .ZN(n2280) );
  AND3_X1 U1758 ( .A1(ADD_RD1[4]), .A2(n2291), .A3(ADD_RD1[0]), .ZN(n2288) );
  AND3_X1 U1759 ( .A1(n2286), .A2(n2291), .A3(ADD_RD1[4]), .ZN(n2289) );
  AND3_X1 U1760 ( .A1(ADD_RD2[4]), .A2(n1659), .A3(ADD_RD2[0]), .ZN(n1654) );
  AND3_X1 U1761 ( .A1(ADD_RD1[4]), .A2(n2286), .A3(ADD_RD1[3]), .ZN(n2281) );
  AND3_X1 U1762 ( .A1(n1650), .A2(n1659), .A3(ADD_RD2[4]), .ZN(n1655) );
  AND3_X1 U1763 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(ADD_RD1[3]), .ZN(n2279) );
  AND3_X1 U1764 ( .A1(ADD_RD2[4]), .A2(n1650), .A3(ADD_RD2[3]), .ZN(n1643) );
  AND3_X1 U1765 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n1641) );
  INV_X1 U1766 ( .A(ADD_RD2[3]), .ZN(n1659) );
  INV_X1 U1767 ( .A(ADD_RD2[0]), .ZN(n1650) );
  INV_X1 U1768 ( .A(ADD_RD1[3]), .ZN(n2291) );
  INV_X1 U1769 ( .A(ADD_RD1[0]), .ZN(n2286) );
  AND2_X1 U1770 ( .A1(WR), .A2(ENABLE), .ZN(n535) );
  BUF_X1 U1771 ( .A(RESET), .Z(n3093) );
  INV_X1 U1772 ( .A(ADD_WR[2]), .ZN(n543) );
  INV_X1 U1773 ( .A(ADD_WR[0]), .ZN(n541) );
  INV_X1 U1774 ( .A(ADD_WR[1]), .ZN(n542) );
  NAND2_X1 U1775 ( .A1(n3097), .A2(n544), .ZN(n2503) );
  NAND2_X1 U1776 ( .A1(RD1), .A2(ENABLE), .ZN(n544) );
  NAND2_X1 U1777 ( .A1(n3097), .A2(n545), .ZN(n2500) );
  NAND2_X1 U1778 ( .A1(RD2), .A2(ENABLE), .ZN(n545) );
  INV_X1 U1779 ( .A(\REGISTERS[28][0] ), .ZN(n1638) );
  INV_X1 U1780 ( .A(\REGISTERS[24][0] ), .ZN(n1645) );
  INV_X1 U1781 ( .A(\REGISTERS[20][0] ), .ZN(n1651) );
  INV_X1 U1782 ( .A(\REGISTERS[16][0] ), .ZN(n1656) );
  INV_X1 U1783 ( .A(\REGISTERS[12][0] ), .ZN(n1664) );
  INV_X1 U1784 ( .A(\REGISTERS[8][0] ), .ZN(n1669) );
  INV_X1 U1785 ( .A(\REGISTERS[4][0] ), .ZN(n1672) );
  INV_X1 U1786 ( .A(\REGISTERS[0][0] ), .ZN(n1678) );
  INV_X1 U1787 ( .A(\REGISTERS[28][1] ), .ZN(n1604) );
  INV_X1 U1788 ( .A(\REGISTERS[24][1] ), .ZN(n1607) );
  INV_X1 U1789 ( .A(\REGISTERS[20][1] ), .ZN(n1610) );
  INV_X1 U1790 ( .A(\REGISTERS[16][1] ), .ZN(n1613) );
  INV_X1 U1791 ( .A(\REGISTERS[12][1] ), .ZN(n1620) );
  INV_X1 U1792 ( .A(\REGISTERS[8][1] ), .ZN(n1623) );
  INV_X1 U1793 ( .A(\REGISTERS[4][1] ), .ZN(n1626) );
  INV_X1 U1794 ( .A(\REGISTERS[0][1] ), .ZN(n1629) );
  INV_X1 U1795 ( .A(\REGISTERS[28][2] ), .ZN(n1570) );
  INV_X1 U1796 ( .A(\REGISTERS[24][2] ), .ZN(n1573) );
  INV_X1 U1797 ( .A(\REGISTERS[20][2] ), .ZN(n1576) );
  INV_X1 U1798 ( .A(\REGISTERS[16][2] ), .ZN(n1579) );
  INV_X1 U1799 ( .A(\REGISTERS[12][2] ), .ZN(n1586) );
  INV_X1 U1800 ( .A(\REGISTERS[8][2] ), .ZN(n1589) );
  INV_X1 U1801 ( .A(\REGISTERS[4][2] ), .ZN(n1592) );
  INV_X1 U1802 ( .A(\REGISTERS[0][2] ), .ZN(n1595) );
  INV_X1 U1803 ( .A(\REGISTERS[28][3] ), .ZN(n1536) );
  INV_X1 U1804 ( .A(\REGISTERS[24][3] ), .ZN(n1539) );
  INV_X1 U1805 ( .A(\REGISTERS[20][3] ), .ZN(n1542) );
  INV_X1 U1806 ( .A(\REGISTERS[16][3] ), .ZN(n1545) );
  INV_X1 U1807 ( .A(\REGISTERS[12][3] ), .ZN(n1552) );
  INV_X1 U1808 ( .A(\REGISTERS[8][3] ), .ZN(n1555) );
  INV_X1 U1809 ( .A(\REGISTERS[4][3] ), .ZN(n1558) );
  INV_X1 U1810 ( .A(\REGISTERS[0][3] ), .ZN(n1561) );
  INV_X1 U1811 ( .A(\REGISTERS[28][4] ), .ZN(n1502) );
  INV_X1 U1812 ( .A(\REGISTERS[24][4] ), .ZN(n1505) );
  INV_X1 U1813 ( .A(\REGISTERS[20][4] ), .ZN(n1508) );
  INV_X1 U1814 ( .A(\REGISTERS[16][4] ), .ZN(n1511) );
  INV_X1 U1815 ( .A(\REGISTERS[12][4] ), .ZN(n1518) );
  INV_X1 U1816 ( .A(\REGISTERS[8][4] ), .ZN(n1521) );
  INV_X1 U1817 ( .A(\REGISTERS[4][4] ), .ZN(n1524) );
  INV_X1 U1818 ( .A(\REGISTERS[0][4] ), .ZN(n1527) );
  INV_X1 U1819 ( .A(\REGISTERS[28][5] ), .ZN(n1468) );
  INV_X1 U1820 ( .A(\REGISTERS[24][5] ), .ZN(n1471) );
  INV_X1 U1821 ( .A(\REGISTERS[20][5] ), .ZN(n1474) );
  INV_X1 U1822 ( .A(\REGISTERS[16][5] ), .ZN(n1477) );
  INV_X1 U1823 ( .A(\REGISTERS[12][5] ), .ZN(n1484) );
  INV_X1 U1824 ( .A(\REGISTERS[8][5] ), .ZN(n1487) );
  INV_X1 U1825 ( .A(\REGISTERS[4][5] ), .ZN(n1490) );
  INV_X1 U1826 ( .A(\REGISTERS[0][5] ), .ZN(n1493) );
  INV_X1 U1827 ( .A(\REGISTERS[28][6] ), .ZN(n1434) );
  INV_X1 U1828 ( .A(\REGISTERS[24][6] ), .ZN(n1437) );
  INV_X1 U1829 ( .A(\REGISTERS[20][6] ), .ZN(n1440) );
  INV_X1 U1830 ( .A(\REGISTERS[16][6] ), .ZN(n1443) );
  INV_X1 U1831 ( .A(\REGISTERS[12][6] ), .ZN(n1450) );
  INV_X1 U1832 ( .A(\REGISTERS[8][6] ), .ZN(n1453) );
  INV_X1 U1833 ( .A(\REGISTERS[4][6] ), .ZN(n1456) );
  INV_X1 U1834 ( .A(\REGISTERS[0][6] ), .ZN(n1459) );
  INV_X1 U1835 ( .A(\REGISTERS[28][7] ), .ZN(n1400) );
  INV_X1 U1836 ( .A(\REGISTERS[24][7] ), .ZN(n1403) );
  INV_X1 U1837 ( .A(\REGISTERS[20][7] ), .ZN(n1406) );
  INV_X1 U1838 ( .A(\REGISTERS[16][7] ), .ZN(n1409) );
  INV_X1 U1839 ( .A(\REGISTERS[12][7] ), .ZN(n1416) );
  INV_X1 U1840 ( .A(\REGISTERS[8][7] ), .ZN(n1419) );
  INV_X1 U1841 ( .A(\REGISTERS[4][7] ), .ZN(n1422) );
  INV_X1 U1842 ( .A(\REGISTERS[0][7] ), .ZN(n1425) );
  INV_X1 U1843 ( .A(\REGISTERS[28][8] ), .ZN(n1366) );
  INV_X1 U1844 ( .A(\REGISTERS[24][8] ), .ZN(n1369) );
  INV_X1 U1845 ( .A(\REGISTERS[20][8] ), .ZN(n1372) );
  INV_X1 U1846 ( .A(\REGISTERS[16][8] ), .ZN(n1375) );
  INV_X1 U1847 ( .A(\REGISTERS[12][8] ), .ZN(n1382) );
  INV_X1 U1848 ( .A(\REGISTERS[8][8] ), .ZN(n1385) );
  INV_X1 U1849 ( .A(\REGISTERS[4][8] ), .ZN(n1388) );
  INV_X1 U1850 ( .A(\REGISTERS[0][8] ), .ZN(n1391) );
  INV_X1 U1851 ( .A(\REGISTERS[28][9] ), .ZN(n1332) );
  INV_X1 U1852 ( .A(\REGISTERS[24][9] ), .ZN(n1335) );
  INV_X1 U1853 ( .A(\REGISTERS[20][9] ), .ZN(n1338) );
  INV_X1 U1854 ( .A(\REGISTERS[16][9] ), .ZN(n1341) );
  INV_X1 U1855 ( .A(\REGISTERS[12][9] ), .ZN(n1348) );
  INV_X1 U1856 ( .A(\REGISTERS[8][9] ), .ZN(n1351) );
  INV_X1 U1857 ( .A(\REGISTERS[4][9] ), .ZN(n1354) );
  INV_X1 U1858 ( .A(\REGISTERS[0][9] ), .ZN(n1357) );
  INV_X1 U1859 ( .A(\REGISTERS[28][10] ), .ZN(n1298) );
  INV_X1 U1860 ( .A(\REGISTERS[24][10] ), .ZN(n1301) );
  INV_X1 U1861 ( .A(\REGISTERS[20][10] ), .ZN(n1304) );
  INV_X1 U1862 ( .A(\REGISTERS[16][10] ), .ZN(n1307) );
  INV_X1 U1863 ( .A(\REGISTERS[12][10] ), .ZN(n1314) );
  INV_X1 U1864 ( .A(\REGISTERS[8][10] ), .ZN(n1317) );
  INV_X1 U1865 ( .A(\REGISTERS[4][10] ), .ZN(n1320) );
  INV_X1 U1866 ( .A(\REGISTERS[0][10] ), .ZN(n1323) );
  INV_X1 U1867 ( .A(\REGISTERS[28][11] ), .ZN(n1264) );
  INV_X1 U1868 ( .A(\REGISTERS[24][11] ), .ZN(n1267) );
  INV_X1 U1869 ( .A(\REGISTERS[20][11] ), .ZN(n1270) );
  INV_X1 U1870 ( .A(\REGISTERS[16][11] ), .ZN(n1273) );
  INV_X1 U1871 ( .A(\REGISTERS[12][11] ), .ZN(n1280) );
  INV_X1 U1872 ( .A(\REGISTERS[8][11] ), .ZN(n1283) );
  INV_X1 U1873 ( .A(\REGISTERS[4][11] ), .ZN(n1286) );
  INV_X1 U1874 ( .A(\REGISTERS[0][11] ), .ZN(n1289) );
  INV_X1 U1875 ( .A(\REGISTERS[28][12] ), .ZN(n1230) );
  INV_X1 U1876 ( .A(\REGISTERS[24][12] ), .ZN(n1233) );
  INV_X1 U1877 ( .A(\REGISTERS[20][12] ), .ZN(n1236) );
  INV_X1 U1878 ( .A(\REGISTERS[16][12] ), .ZN(n1239) );
  INV_X1 U1879 ( .A(\REGISTERS[12][12] ), .ZN(n1246) );
  INV_X1 U1880 ( .A(\REGISTERS[8][12] ), .ZN(n1249) );
  INV_X1 U1881 ( .A(\REGISTERS[4][12] ), .ZN(n1252) );
  INV_X1 U1882 ( .A(\REGISTERS[0][12] ), .ZN(n1255) );
  INV_X1 U1883 ( .A(\REGISTERS[28][13] ), .ZN(n1196) );
  INV_X1 U1884 ( .A(\REGISTERS[24][13] ), .ZN(n1199) );
  INV_X1 U1885 ( .A(\REGISTERS[20][13] ), .ZN(n1202) );
  INV_X1 U1886 ( .A(\REGISTERS[16][13] ), .ZN(n1205) );
  INV_X1 U1887 ( .A(\REGISTERS[12][13] ), .ZN(n1212) );
  INV_X1 U1888 ( .A(\REGISTERS[8][13] ), .ZN(n1215) );
  INV_X1 U1889 ( .A(\REGISTERS[4][13] ), .ZN(n1218) );
  INV_X1 U1890 ( .A(\REGISTERS[0][13] ), .ZN(n1221) );
  INV_X1 U1891 ( .A(\REGISTERS[28][14] ), .ZN(n1162) );
  INV_X1 U1892 ( .A(\REGISTERS[24][14] ), .ZN(n1165) );
  INV_X1 U1893 ( .A(\REGISTERS[20][14] ), .ZN(n1168) );
  INV_X1 U1894 ( .A(\REGISTERS[16][14] ), .ZN(n1171) );
  INV_X1 U1895 ( .A(\REGISTERS[12][14] ), .ZN(n1178) );
  INV_X1 U1896 ( .A(\REGISTERS[8][14] ), .ZN(n1181) );
  INV_X1 U1897 ( .A(\REGISTERS[4][14] ), .ZN(n1184) );
  INV_X1 U1898 ( .A(\REGISTERS[0][14] ), .ZN(n1187) );
  INV_X1 U1899 ( .A(\REGISTERS[28][15] ), .ZN(n1128) );
  INV_X1 U1900 ( .A(\REGISTERS[24][15] ), .ZN(n1131) );
  INV_X1 U1913 ( .A(\REGISTERS[20][15] ), .ZN(n1134) );
  INV_X1 U1914 ( .A(\REGISTERS[16][15] ), .ZN(n1137) );
  INV_X1 U1915 ( .A(\REGISTERS[12][15] ), .ZN(n1144) );
  INV_X1 U1916 ( .A(\REGISTERS[8][15] ), .ZN(n1147) );
  INV_X1 U1917 ( .A(\REGISTERS[4][15] ), .ZN(n1150) );
  INV_X1 U1918 ( .A(\REGISTERS[0][15] ), .ZN(n1153) );
  INV_X1 U1919 ( .A(\REGISTERS[28][16] ), .ZN(n1094) );
  INV_X1 U1920 ( .A(\REGISTERS[24][16] ), .ZN(n1097) );
  INV_X1 U1921 ( .A(\REGISTERS[20][16] ), .ZN(n1100) );
  INV_X1 U1922 ( .A(\REGISTERS[16][16] ), .ZN(n1103) );
  INV_X1 U1923 ( .A(\REGISTERS[12][16] ), .ZN(n1110) );
  INV_X1 U1924 ( .A(\REGISTERS[8][16] ), .ZN(n1113) );
  INV_X1 U1925 ( .A(\REGISTERS[4][16] ), .ZN(n1116) );
  INV_X1 U1926 ( .A(\REGISTERS[0][16] ), .ZN(n1119) );
  INV_X1 U1927 ( .A(\REGISTERS[28][17] ), .ZN(n1060) );
  INV_X1 U1928 ( .A(\REGISTERS[24][17] ), .ZN(n1063) );
  INV_X1 U1929 ( .A(\REGISTERS[20][17] ), .ZN(n1066) );
  INV_X1 U1930 ( .A(\REGISTERS[16][17] ), .ZN(n1069) );
  INV_X1 U1931 ( .A(\REGISTERS[12][17] ), .ZN(n1076) );
  INV_X1 U1932 ( .A(\REGISTERS[8][17] ), .ZN(n1079) );
  INV_X1 U1933 ( .A(\REGISTERS[4][17] ), .ZN(n1082) );
  INV_X1 U1934 ( .A(\REGISTERS[0][17] ), .ZN(n1085) );
  INV_X1 U1935 ( .A(\REGISTERS[28][18] ), .ZN(n1026) );
  INV_X1 U1936 ( .A(\REGISTERS[24][18] ), .ZN(n1029) );
  INV_X1 U1937 ( .A(\REGISTERS[20][18] ), .ZN(n1032) );
  INV_X1 U1938 ( .A(\REGISTERS[16][18] ), .ZN(n1035) );
  INV_X1 U1939 ( .A(\REGISTERS[12][18] ), .ZN(n1042) );
  INV_X1 U1940 ( .A(\REGISTERS[8][18] ), .ZN(n1045) );
  INV_X1 U1941 ( .A(\REGISTERS[4][18] ), .ZN(n1048) );
  INV_X1 U1942 ( .A(\REGISTERS[0][18] ), .ZN(n1051) );
  INV_X1 U1943 ( .A(\REGISTERS[28][19] ), .ZN(n992) );
  INV_X1 U1944 ( .A(\REGISTERS[24][19] ), .ZN(n995) );
  INV_X1 U1945 ( .A(\REGISTERS[20][19] ), .ZN(n998) );
  INV_X1 U1946 ( .A(\REGISTERS[16][19] ), .ZN(n1001) );
  INV_X1 U1947 ( .A(\REGISTERS[12][19] ), .ZN(n1008) );
  INV_X1 U1948 ( .A(\REGISTERS[8][19] ), .ZN(n1011) );
  INV_X1 U1949 ( .A(\REGISTERS[4][19] ), .ZN(n1014) );
  INV_X1 U1950 ( .A(\REGISTERS[0][19] ), .ZN(n1017) );
  INV_X1 U1951 ( .A(\REGISTERS[28][20] ), .ZN(n958) );
  INV_X1 U1952 ( .A(\REGISTERS[24][20] ), .ZN(n961) );
  INV_X1 U1953 ( .A(\REGISTERS[20][20] ), .ZN(n964) );
  INV_X1 U1954 ( .A(\REGISTERS[16][20] ), .ZN(n967) );
  INV_X1 U1955 ( .A(\REGISTERS[12][20] ), .ZN(n974) );
  INV_X1 U1956 ( .A(\REGISTERS[8][20] ), .ZN(n977) );
  INV_X1 U1957 ( .A(\REGISTERS[4][20] ), .ZN(n980) );
  INV_X1 U1958 ( .A(\REGISTERS[0][20] ), .ZN(n983) );
  INV_X1 U1959 ( .A(\REGISTERS[28][21] ), .ZN(n924) );
  INV_X1 U1960 ( .A(\REGISTERS[24][21] ), .ZN(n927) );
  INV_X1 U1961 ( .A(\REGISTERS[20][21] ), .ZN(n930) );
  INV_X1 U1962 ( .A(\REGISTERS[16][21] ), .ZN(n933) );
  INV_X1 U1963 ( .A(\REGISTERS[12][21] ), .ZN(n940) );
  INV_X1 U1964 ( .A(\REGISTERS[8][21] ), .ZN(n943) );
  INV_X1 U1965 ( .A(\REGISTERS[4][21] ), .ZN(n946) );
  INV_X1 U1966 ( .A(\REGISTERS[0][21] ), .ZN(n949) );
  INV_X1 U1967 ( .A(\REGISTERS[28][22] ), .ZN(n890) );
  INV_X1 U1968 ( .A(\REGISTERS[24][22] ), .ZN(n893) );
  INV_X1 U1969 ( .A(\REGISTERS[20][22] ), .ZN(n896) );
  INV_X1 U1970 ( .A(\REGISTERS[16][22] ), .ZN(n899) );
  INV_X1 U1971 ( .A(\REGISTERS[12][22] ), .ZN(n906) );
  INV_X1 U1972 ( .A(\REGISTERS[8][22] ), .ZN(n909) );
  INV_X1 U1973 ( .A(\REGISTERS[4][22] ), .ZN(n912) );
  INV_X1 U1974 ( .A(\REGISTERS[0][22] ), .ZN(n915) );
  INV_X1 U1975 ( .A(\REGISTERS[28][23] ), .ZN(n856) );
  INV_X1 U1976 ( .A(\REGISTERS[24][23] ), .ZN(n859) );
  INV_X1 U1977 ( .A(\REGISTERS[20][23] ), .ZN(n862) );
  INV_X1 U1978 ( .A(\REGISTERS[16][23] ), .ZN(n865) );
  INV_X1 U1979 ( .A(\REGISTERS[12][23] ), .ZN(n872) );
  INV_X1 U1980 ( .A(\REGISTERS[8][23] ), .ZN(n875) );
  INV_X1 U1981 ( .A(\REGISTERS[4][23] ), .ZN(n878) );
  INV_X1 U1982 ( .A(\REGISTERS[0][23] ), .ZN(n881) );
  INV_X1 U1983 ( .A(\REGISTERS[28][24] ), .ZN(n822) );
  INV_X1 U1984 ( .A(\REGISTERS[24][24] ), .ZN(n825) );
  INV_X1 U1985 ( .A(\REGISTERS[20][24] ), .ZN(n828) );
  INV_X1 U1986 ( .A(\REGISTERS[16][24] ), .ZN(n831) );
  INV_X1 U1987 ( .A(\REGISTERS[12][24] ), .ZN(n838) );
  INV_X1 U1988 ( .A(\REGISTERS[8][24] ), .ZN(n841) );
  INV_X1 U1989 ( .A(\REGISTERS[4][24] ), .ZN(n844) );
  INV_X1 U1990 ( .A(\REGISTERS[0][24] ), .ZN(n847) );
  INV_X1 U1991 ( .A(\REGISTERS[28][25] ), .ZN(n788) );
  INV_X1 U1992 ( .A(\REGISTERS[24][25] ), .ZN(n791) );
  INV_X1 U1993 ( .A(\REGISTERS[20][25] ), .ZN(n794) );
  INV_X1 U1994 ( .A(\REGISTERS[16][25] ), .ZN(n797) );
  INV_X1 U1995 ( .A(\REGISTERS[12][25] ), .ZN(n804) );
  INV_X1 U1996 ( .A(\REGISTERS[8][25] ), .ZN(n807) );
  INV_X1 U1997 ( .A(\REGISTERS[4][25] ), .ZN(n810) );
  INV_X1 U1998 ( .A(\REGISTERS[0][25] ), .ZN(n813) );
  INV_X1 U1999 ( .A(\REGISTERS[28][26] ), .ZN(n754) );
  INV_X1 U2000 ( .A(\REGISTERS[24][26] ), .ZN(n757) );
  INV_X1 U2001 ( .A(\REGISTERS[20][26] ), .ZN(n760) );
  INV_X1 U2002 ( .A(\REGISTERS[16][26] ), .ZN(n763) );
  INV_X1 U2003 ( .A(\REGISTERS[12][26] ), .ZN(n770) );
  INV_X1 U2004 ( .A(\REGISTERS[8][26] ), .ZN(n773) );
  INV_X1 U2005 ( .A(\REGISTERS[4][26] ), .ZN(n776) );
  INV_X1 U2006 ( .A(\REGISTERS[0][26] ), .ZN(n779) );
  INV_X1 U2007 ( .A(\REGISTERS[28][27] ), .ZN(n720) );
  INV_X1 U2008 ( .A(\REGISTERS[24][27] ), .ZN(n723) );
  INV_X1 U2009 ( .A(\REGISTERS[20][27] ), .ZN(n726) );
  INV_X1 U2010 ( .A(\REGISTERS[16][27] ), .ZN(n729) );
  INV_X1 U2011 ( .A(\REGISTERS[12][27] ), .ZN(n736) );
  INV_X1 U2012 ( .A(\REGISTERS[8][27] ), .ZN(n739) );
  INV_X1 U2013 ( .A(\REGISTERS[4][27] ), .ZN(n742) );
  INV_X1 U2014 ( .A(\REGISTERS[0][27] ), .ZN(n745) );
  INV_X1 U2015 ( .A(\REGISTERS[28][28] ), .ZN(n686) );
  INV_X1 U2016 ( .A(\REGISTERS[24][28] ), .ZN(n689) );
  INV_X1 U2017 ( .A(\REGISTERS[20][28] ), .ZN(n692) );
  INV_X1 U2018 ( .A(\REGISTERS[16][28] ), .ZN(n695) );
  INV_X1 U2019 ( .A(\REGISTERS[12][28] ), .ZN(n702) );
  INV_X1 U2020 ( .A(\REGISTERS[8][28] ), .ZN(n705) );
  INV_X1 U2021 ( .A(\REGISTERS[4][28] ), .ZN(n708) );
  INV_X1 U2022 ( .A(\REGISTERS[0][28] ), .ZN(n711) );
  INV_X1 U2023 ( .A(\REGISTERS[28][29] ), .ZN(n652) );
  INV_X1 U2024 ( .A(\REGISTERS[24][29] ), .ZN(n655) );
  INV_X1 U2025 ( .A(\REGISTERS[20][29] ), .ZN(n658) );
  INV_X1 U2026 ( .A(\REGISTERS[16][29] ), .ZN(n661) );
  INV_X1 U2027 ( .A(\REGISTERS[12][29] ), .ZN(n668) );
  INV_X1 U2028 ( .A(\REGISTERS[8][29] ), .ZN(n671) );
  INV_X1 U2029 ( .A(\REGISTERS[4][29] ), .ZN(n674) );
  INV_X1 U2030 ( .A(\REGISTERS[0][29] ), .ZN(n677) );
  INV_X1 U2031 ( .A(\REGISTERS[28][30] ), .ZN(n618) );
  INV_X1 U2032 ( .A(\REGISTERS[24][30] ), .ZN(n621) );
  INV_X1 U2033 ( .A(\REGISTERS[20][30] ), .ZN(n624) );
  INV_X1 U2034 ( .A(\REGISTERS[16][30] ), .ZN(n627) );
  INV_X1 U2035 ( .A(\REGISTERS[12][30] ), .ZN(n634) );
  INV_X1 U2036 ( .A(\REGISTERS[8][30] ), .ZN(n637) );
  INV_X1 U2037 ( .A(\REGISTERS[4][30] ), .ZN(n640) );
  INV_X1 U2038 ( .A(\REGISTERS[0][30] ), .ZN(n643) );
  INV_X1 U2039 ( .A(\REGISTERS[28][31] ), .ZN(n553) );
  INV_X1 U2040 ( .A(\REGISTERS[24][31] ), .ZN(n560) );
  INV_X1 U2041 ( .A(\REGISTERS[20][31] ), .ZN(n567) );
  INV_X1 U2042 ( .A(\REGISTERS[16][31] ), .ZN(n574) );
  INV_X1 U2043 ( .A(\REGISTERS[12][31] ), .ZN(n585) );
  INV_X1 U2044 ( .A(\REGISTERS[8][31] ), .ZN(n592) );
  INV_X1 U2045 ( .A(\REGISTERS[4][31] ), .ZN(n599) );
  INV_X1 U2046 ( .A(\REGISTERS[0][31] ), .ZN(n606) );
  INV_X1 U2047 ( .A(\REGISTERS[29][0] ), .ZN(n1639) );
  INV_X1 U2048 ( .A(\REGISTERS[25][0] ), .ZN(n1646) );
  INV_X1 U2049 ( .A(\REGISTERS[21][0] ), .ZN(n1652) );
  INV_X1 U2050 ( .A(\REGISTERS[17][0] ), .ZN(n1657) );
  INV_X1 U2051 ( .A(\REGISTERS[13][0] ), .ZN(n1665) );
  INV_X1 U2052 ( .A(\REGISTERS[9][0] ), .ZN(n1670) );
  INV_X1 U2053 ( .A(\REGISTERS[5][0] ), .ZN(n1673) );
  INV_X1 U2054 ( .A(\REGISTERS[1][0] ), .ZN(n1679) );
  INV_X1 U2055 ( .A(\REGISTERS[29][1] ), .ZN(n1605) );
  INV_X1 U2056 ( .A(\REGISTERS[25][1] ), .ZN(n1608) );
  INV_X1 U2057 ( .A(\REGISTERS[21][1] ), .ZN(n1611) );
  INV_X1 U2058 ( .A(\REGISTERS[17][1] ), .ZN(n1614) );
  INV_X1 U2059 ( .A(\REGISTERS[13][1] ), .ZN(n1621) );
  INV_X1 U2060 ( .A(\REGISTERS[9][1] ), .ZN(n1624) );
  INV_X1 U2061 ( .A(\REGISTERS[5][1] ), .ZN(n1627) );
  INV_X1 U2062 ( .A(\REGISTERS[1][1] ), .ZN(n1630) );
  INV_X1 U2063 ( .A(\REGISTERS[29][2] ), .ZN(n1571) );
  INV_X1 U2064 ( .A(\REGISTERS[25][2] ), .ZN(n1574) );
  INV_X1 U2065 ( .A(\REGISTERS[21][2] ), .ZN(n1577) );
  INV_X1 U2066 ( .A(\REGISTERS[17][2] ), .ZN(n1580) );
  INV_X1 U2067 ( .A(\REGISTERS[13][2] ), .ZN(n1587) );
  INV_X1 U2068 ( .A(\REGISTERS[9][2] ), .ZN(n1590) );
  INV_X1 U2069 ( .A(\REGISTERS[5][2] ), .ZN(n1593) );
  INV_X1 U2070 ( .A(\REGISTERS[1][2] ), .ZN(n1596) );
  INV_X1 U2071 ( .A(\REGISTERS[29][3] ), .ZN(n1537) );
  INV_X1 U2072 ( .A(\REGISTERS[25][3] ), .ZN(n1540) );
  INV_X1 U2073 ( .A(\REGISTERS[21][3] ), .ZN(n1543) );
  INV_X1 U2074 ( .A(\REGISTERS[17][3] ), .ZN(n1546) );
  INV_X1 U2075 ( .A(\REGISTERS[13][3] ), .ZN(n1553) );
  INV_X1 U2076 ( .A(\REGISTERS[9][3] ), .ZN(n1556) );
  INV_X1 U2077 ( .A(\REGISTERS[5][3] ), .ZN(n1559) );
  INV_X1 U2078 ( .A(\REGISTERS[1][3] ), .ZN(n1562) );
  INV_X1 U2079 ( .A(\REGISTERS[29][4] ), .ZN(n1503) );
  INV_X1 U2080 ( .A(\REGISTERS[25][4] ), .ZN(n1506) );
  INV_X1 U2081 ( .A(\REGISTERS[21][4] ), .ZN(n1509) );
  INV_X1 U2082 ( .A(\REGISTERS[17][4] ), .ZN(n1512) );
  INV_X1 U2083 ( .A(\REGISTERS[13][4] ), .ZN(n1519) );
  INV_X1 U2084 ( .A(\REGISTERS[9][4] ), .ZN(n1522) );
  INV_X1 U2085 ( .A(\REGISTERS[5][4] ), .ZN(n1525) );
  INV_X1 U2086 ( .A(\REGISTERS[1][4] ), .ZN(n1528) );
  INV_X1 U2087 ( .A(\REGISTERS[29][5] ), .ZN(n1469) );
  INV_X1 U2088 ( .A(\REGISTERS[25][5] ), .ZN(n1472) );
  INV_X1 U2089 ( .A(\REGISTERS[21][5] ), .ZN(n1475) );
  INV_X1 U2090 ( .A(\REGISTERS[17][5] ), .ZN(n1478) );
  INV_X1 U2091 ( .A(\REGISTERS[13][5] ), .ZN(n1485) );
  INV_X1 U2092 ( .A(\REGISTERS[9][5] ), .ZN(n1488) );
  INV_X1 U2093 ( .A(\REGISTERS[5][5] ), .ZN(n1491) );
  INV_X1 U2094 ( .A(\REGISTERS[1][5] ), .ZN(n1494) );
  INV_X1 U2095 ( .A(\REGISTERS[29][6] ), .ZN(n1435) );
  INV_X1 U2096 ( .A(\REGISTERS[25][6] ), .ZN(n1438) );
  INV_X1 U2097 ( .A(\REGISTERS[21][6] ), .ZN(n1441) );
  INV_X1 U2098 ( .A(\REGISTERS[17][6] ), .ZN(n1444) );
  INV_X1 U2099 ( .A(\REGISTERS[13][6] ), .ZN(n1451) );
  INV_X1 U2100 ( .A(\REGISTERS[9][6] ), .ZN(n1454) );
  INV_X1 U2101 ( .A(\REGISTERS[5][6] ), .ZN(n1457) );
  INV_X1 U2102 ( .A(\REGISTERS[1][6] ), .ZN(n1460) );
  INV_X1 U2103 ( .A(\REGISTERS[29][7] ), .ZN(n1401) );
  INV_X1 U2104 ( .A(\REGISTERS[25][7] ), .ZN(n1404) );
  INV_X1 U2105 ( .A(\REGISTERS[21][7] ), .ZN(n1407) );
  INV_X1 U2106 ( .A(\REGISTERS[17][7] ), .ZN(n1410) );
  INV_X1 U2107 ( .A(\REGISTERS[13][7] ), .ZN(n1417) );
  INV_X1 U2108 ( .A(\REGISTERS[9][7] ), .ZN(n1420) );
  INV_X1 U2109 ( .A(\REGISTERS[5][7] ), .ZN(n1423) );
  INV_X1 U2110 ( .A(\REGISTERS[1][7] ), .ZN(n1426) );
  INV_X1 U2111 ( .A(\REGISTERS[29][8] ), .ZN(n1367) );
  INV_X1 U2112 ( .A(\REGISTERS[25][8] ), .ZN(n1370) );
  INV_X1 U2113 ( .A(\REGISTERS[21][8] ), .ZN(n1373) );
  INV_X1 U2114 ( .A(\REGISTERS[17][8] ), .ZN(n1376) );
  INV_X1 U2115 ( .A(\REGISTERS[13][8] ), .ZN(n1383) );
  INV_X1 U2116 ( .A(\REGISTERS[9][8] ), .ZN(n1386) );
  INV_X1 U2117 ( .A(\REGISTERS[5][8] ), .ZN(n1389) );
  INV_X1 U2118 ( .A(\REGISTERS[1][8] ), .ZN(n1392) );
  INV_X1 U2119 ( .A(\REGISTERS[29][9] ), .ZN(n1333) );
  INV_X1 U2120 ( .A(\REGISTERS[25][9] ), .ZN(n1336) );
  INV_X1 U2121 ( .A(\REGISTERS[21][9] ), .ZN(n1339) );
  INV_X1 U2122 ( .A(\REGISTERS[17][9] ), .ZN(n1342) );
  INV_X1 U2123 ( .A(\REGISTERS[13][9] ), .ZN(n1349) );
  INV_X1 U2124 ( .A(\REGISTERS[9][9] ), .ZN(n1352) );
  INV_X1 U2125 ( .A(\REGISTERS[5][9] ), .ZN(n1355) );
  INV_X1 U2126 ( .A(\REGISTERS[1][9] ), .ZN(n1358) );
  INV_X1 U2127 ( .A(\REGISTERS[29][10] ), .ZN(n1299) );
  INV_X1 U2128 ( .A(\REGISTERS[25][10] ), .ZN(n1302) );
  INV_X1 U2129 ( .A(\REGISTERS[21][10] ), .ZN(n1305) );
  INV_X1 U2130 ( .A(\REGISTERS[17][10] ), .ZN(n1308) );
  INV_X1 U2131 ( .A(\REGISTERS[13][10] ), .ZN(n1315) );
  INV_X1 U2132 ( .A(\REGISTERS[9][10] ), .ZN(n1318) );
  INV_X1 U2133 ( .A(\REGISTERS[5][10] ), .ZN(n1321) );
  INV_X1 U2134 ( .A(\REGISTERS[1][10] ), .ZN(n1324) );
  INV_X1 U2135 ( .A(\REGISTERS[29][11] ), .ZN(n1265) );
  INV_X1 U2136 ( .A(\REGISTERS[25][11] ), .ZN(n1268) );
  INV_X1 U2137 ( .A(\REGISTERS[21][11] ), .ZN(n1271) );
  INV_X1 U2138 ( .A(\REGISTERS[17][11] ), .ZN(n1274) );
  INV_X1 U2139 ( .A(\REGISTERS[13][11] ), .ZN(n1281) );
  INV_X1 U2140 ( .A(\REGISTERS[9][11] ), .ZN(n1284) );
  INV_X1 U2141 ( .A(\REGISTERS[5][11] ), .ZN(n1287) );
  INV_X1 U2142 ( .A(\REGISTERS[1][11] ), .ZN(n1290) );
  INV_X1 U2143 ( .A(\REGISTERS[29][12] ), .ZN(n1231) );
  INV_X1 U2144 ( .A(\REGISTERS[25][12] ), .ZN(n1234) );
  INV_X1 U2145 ( .A(\REGISTERS[21][12] ), .ZN(n1237) );
  INV_X1 U2146 ( .A(\REGISTERS[17][12] ), .ZN(n1240) );
  INV_X1 U2147 ( .A(\REGISTERS[13][12] ), .ZN(n1247) );
  INV_X1 U2148 ( .A(\REGISTERS[9][12] ), .ZN(n1250) );
  INV_X1 U2149 ( .A(\REGISTERS[5][12] ), .ZN(n1253) );
  INV_X1 U2150 ( .A(\REGISTERS[1][12] ), .ZN(n1256) );
  INV_X1 U2151 ( .A(\REGISTERS[29][13] ), .ZN(n1197) );
  INV_X1 U2152 ( .A(\REGISTERS[25][13] ), .ZN(n1200) );
  INV_X1 U2153 ( .A(\REGISTERS[21][13] ), .ZN(n1203) );
  INV_X1 U2154 ( .A(\REGISTERS[17][13] ), .ZN(n1206) );
  INV_X1 U2155 ( .A(\REGISTERS[13][13] ), .ZN(n1213) );
  INV_X1 U2156 ( .A(\REGISTERS[9][13] ), .ZN(n1216) );
  INV_X1 U2157 ( .A(\REGISTERS[5][13] ), .ZN(n1219) );
  INV_X1 U2158 ( .A(\REGISTERS[1][13] ), .ZN(n1222) );
  INV_X1 U2159 ( .A(\REGISTERS[29][14] ), .ZN(n1163) );
  INV_X1 U2160 ( .A(\REGISTERS[25][14] ), .ZN(n1166) );
  INV_X1 U2161 ( .A(\REGISTERS[21][14] ), .ZN(n1169) );
  INV_X1 U2162 ( .A(\REGISTERS[17][14] ), .ZN(n1172) );
  INV_X1 U2163 ( .A(\REGISTERS[13][14] ), .ZN(n1179) );
  INV_X1 U2164 ( .A(\REGISTERS[9][14] ), .ZN(n1182) );
  INV_X1 U2165 ( .A(\REGISTERS[5][14] ), .ZN(n1185) );
  INV_X1 U2166 ( .A(\REGISTERS[1][14] ), .ZN(n1188) );
  INV_X1 U2167 ( .A(\REGISTERS[29][15] ), .ZN(n1129) );
  INV_X1 U2168 ( .A(\REGISTERS[25][15] ), .ZN(n1132) );
  INV_X1 U2169 ( .A(\REGISTERS[21][15] ), .ZN(n1135) );
  INV_X1 U2170 ( .A(\REGISTERS[17][15] ), .ZN(n1138) );
  INV_X1 U2171 ( .A(\REGISTERS[13][15] ), .ZN(n1145) );
  INV_X1 U2172 ( .A(\REGISTERS[9][15] ), .ZN(n1148) );
  INV_X1 U2173 ( .A(\REGISTERS[5][15] ), .ZN(n1151) );
  INV_X1 U2174 ( .A(\REGISTERS[1][15] ), .ZN(n1154) );
  INV_X1 U2175 ( .A(\REGISTERS[29][16] ), .ZN(n1095) );
  INV_X1 U2176 ( .A(\REGISTERS[25][16] ), .ZN(n1098) );
  INV_X1 U2177 ( .A(\REGISTERS[21][16] ), .ZN(n1101) );
  INV_X1 U2178 ( .A(\REGISTERS[17][16] ), .ZN(n1104) );
  INV_X1 U2179 ( .A(\REGISTERS[13][16] ), .ZN(n1111) );
  INV_X1 U2180 ( .A(\REGISTERS[9][16] ), .ZN(n1114) );
  INV_X1 U2181 ( .A(\REGISTERS[5][16] ), .ZN(n1117) );
  INV_X1 U2182 ( .A(\REGISTERS[1][16] ), .ZN(n1120) );
  INV_X1 U2183 ( .A(\REGISTERS[29][17] ), .ZN(n1061) );
  INV_X1 U2184 ( .A(\REGISTERS[25][17] ), .ZN(n1064) );
  INV_X1 U2185 ( .A(\REGISTERS[21][17] ), .ZN(n1067) );
  INV_X1 U2186 ( .A(\REGISTERS[17][17] ), .ZN(n1070) );
  INV_X1 U2187 ( .A(\REGISTERS[13][17] ), .ZN(n1077) );
  INV_X1 U2188 ( .A(\REGISTERS[9][17] ), .ZN(n1080) );
  INV_X1 U2189 ( .A(\REGISTERS[5][17] ), .ZN(n1083) );
  INV_X1 U2190 ( .A(\REGISTERS[1][17] ), .ZN(n1086) );
  INV_X1 U2191 ( .A(\REGISTERS[29][18] ), .ZN(n1027) );
  INV_X1 U2192 ( .A(\REGISTERS[25][18] ), .ZN(n1030) );
  INV_X1 U2193 ( .A(\REGISTERS[21][18] ), .ZN(n1033) );
  INV_X1 U2194 ( .A(\REGISTERS[17][18] ), .ZN(n1036) );
  INV_X1 U2195 ( .A(\REGISTERS[13][18] ), .ZN(n1043) );
  INV_X1 U2196 ( .A(\REGISTERS[9][18] ), .ZN(n1046) );
  INV_X1 U2197 ( .A(\REGISTERS[5][18] ), .ZN(n1049) );
  INV_X1 U2198 ( .A(\REGISTERS[1][18] ), .ZN(n1052) );
  INV_X1 U2199 ( .A(\REGISTERS[29][19] ), .ZN(n993) );
  INV_X1 U2200 ( .A(\REGISTERS[25][19] ), .ZN(n996) );
  INV_X1 U2201 ( .A(\REGISTERS[21][19] ), .ZN(n999) );
  INV_X1 U2202 ( .A(\REGISTERS[17][19] ), .ZN(n1002) );
  INV_X1 U2203 ( .A(\REGISTERS[13][19] ), .ZN(n1009) );
  INV_X1 U2204 ( .A(\REGISTERS[9][19] ), .ZN(n1012) );
  INV_X1 U2205 ( .A(\REGISTERS[5][19] ), .ZN(n1015) );
  INV_X1 U2206 ( .A(\REGISTERS[1][19] ), .ZN(n1018) );
  INV_X1 U2207 ( .A(\REGISTERS[29][20] ), .ZN(n959) );
  INV_X1 U2208 ( .A(\REGISTERS[25][20] ), .ZN(n962) );
  INV_X1 U2209 ( .A(\REGISTERS[21][20] ), .ZN(n965) );
  INV_X1 U2210 ( .A(\REGISTERS[17][20] ), .ZN(n968) );
  INV_X1 U2211 ( .A(\REGISTERS[13][20] ), .ZN(n975) );
  INV_X1 U2212 ( .A(\REGISTERS[9][20] ), .ZN(n978) );
  INV_X1 U2213 ( .A(\REGISTERS[5][20] ), .ZN(n981) );
  INV_X1 U2214 ( .A(\REGISTERS[1][20] ), .ZN(n984) );
  INV_X1 U2215 ( .A(\REGISTERS[29][21] ), .ZN(n925) );
  INV_X1 U2216 ( .A(\REGISTERS[25][21] ), .ZN(n928) );
  INV_X1 U2217 ( .A(\REGISTERS[21][21] ), .ZN(n931) );
  INV_X1 U2218 ( .A(\REGISTERS[17][21] ), .ZN(n934) );
  INV_X1 U2219 ( .A(\REGISTERS[13][21] ), .ZN(n941) );
  INV_X1 U2220 ( .A(\REGISTERS[9][21] ), .ZN(n944) );
  INV_X1 U2221 ( .A(\REGISTERS[5][21] ), .ZN(n947) );
  INV_X1 U2222 ( .A(\REGISTERS[1][21] ), .ZN(n950) );
  INV_X1 U2223 ( .A(\REGISTERS[29][22] ), .ZN(n891) );
  INV_X1 U2224 ( .A(\REGISTERS[25][22] ), .ZN(n894) );
  INV_X1 U2225 ( .A(\REGISTERS[21][22] ), .ZN(n897) );
  INV_X1 U2226 ( .A(\REGISTERS[17][22] ), .ZN(n900) );
  INV_X1 U2227 ( .A(\REGISTERS[13][22] ), .ZN(n907) );
  INV_X1 U2228 ( .A(\REGISTERS[9][22] ), .ZN(n910) );
  INV_X1 U2229 ( .A(\REGISTERS[5][22] ), .ZN(n913) );
  INV_X1 U2230 ( .A(\REGISTERS[1][22] ), .ZN(n916) );
  INV_X1 U2231 ( .A(\REGISTERS[29][23] ), .ZN(n857) );
  INV_X1 U2232 ( .A(\REGISTERS[25][23] ), .ZN(n860) );
  INV_X1 U2233 ( .A(\REGISTERS[21][23] ), .ZN(n863) );
  INV_X1 U2234 ( .A(\REGISTERS[17][23] ), .ZN(n866) );
  INV_X1 U2235 ( .A(\REGISTERS[13][23] ), .ZN(n873) );
  INV_X1 U2236 ( .A(\REGISTERS[9][23] ), .ZN(n876) );
  INV_X1 U2237 ( .A(\REGISTERS[5][23] ), .ZN(n879) );
  INV_X1 U2238 ( .A(\REGISTERS[1][23] ), .ZN(n882) );
  INV_X1 U2239 ( .A(\REGISTERS[29][24] ), .ZN(n823) );
  INV_X1 U2240 ( .A(\REGISTERS[25][24] ), .ZN(n826) );
  INV_X1 U2241 ( .A(\REGISTERS[21][24] ), .ZN(n829) );
  INV_X1 U2242 ( .A(\REGISTERS[17][24] ), .ZN(n832) );
  INV_X1 U2243 ( .A(\REGISTERS[13][24] ), .ZN(n839) );
  INV_X1 U2244 ( .A(\REGISTERS[9][24] ), .ZN(n842) );
  INV_X1 U2245 ( .A(\REGISTERS[5][24] ), .ZN(n845) );
  INV_X1 U2246 ( .A(\REGISTERS[1][24] ), .ZN(n848) );
  INV_X1 U2247 ( .A(\REGISTERS[29][25] ), .ZN(n789) );
  INV_X1 U2248 ( .A(\REGISTERS[25][25] ), .ZN(n792) );
  INV_X1 U2249 ( .A(\REGISTERS[21][25] ), .ZN(n795) );
  INV_X1 U2250 ( .A(\REGISTERS[17][25] ), .ZN(n798) );
  INV_X1 U2251 ( .A(\REGISTERS[13][25] ), .ZN(n805) );
  INV_X1 U2252 ( .A(\REGISTERS[9][25] ), .ZN(n808) );
  INV_X1 U2253 ( .A(\REGISTERS[5][25] ), .ZN(n811) );
  INV_X1 U2254 ( .A(\REGISTERS[1][25] ), .ZN(n814) );
  INV_X1 U2255 ( .A(\REGISTERS[29][26] ), .ZN(n755) );
  INV_X1 U2256 ( .A(\REGISTERS[25][26] ), .ZN(n758) );
  INV_X1 U2257 ( .A(\REGISTERS[21][26] ), .ZN(n761) );
  INV_X1 U2258 ( .A(\REGISTERS[17][26] ), .ZN(n764) );
  INV_X1 U2259 ( .A(\REGISTERS[13][26] ), .ZN(n771) );
  INV_X1 U2260 ( .A(\REGISTERS[9][26] ), .ZN(n774) );
  INV_X1 U2261 ( .A(\REGISTERS[5][26] ), .ZN(n777) );
  INV_X1 U2262 ( .A(\REGISTERS[1][26] ), .ZN(n780) );
  INV_X1 U2263 ( .A(\REGISTERS[29][27] ), .ZN(n721) );
  INV_X1 U2264 ( .A(\REGISTERS[25][27] ), .ZN(n724) );
  INV_X1 U2265 ( .A(\REGISTERS[21][27] ), .ZN(n727) );
  INV_X1 U2266 ( .A(\REGISTERS[17][27] ), .ZN(n730) );
  INV_X1 U2267 ( .A(\REGISTERS[13][27] ), .ZN(n737) );
  INV_X1 U2268 ( .A(\REGISTERS[9][27] ), .ZN(n740) );
  INV_X1 U2269 ( .A(\REGISTERS[5][27] ), .ZN(n743) );
  INV_X1 U2270 ( .A(\REGISTERS[1][27] ), .ZN(n746) );
  INV_X1 U2271 ( .A(\REGISTERS[29][28] ), .ZN(n687) );
  INV_X1 U2272 ( .A(\REGISTERS[25][28] ), .ZN(n690) );
  INV_X1 U2273 ( .A(\REGISTERS[21][28] ), .ZN(n693) );
  INV_X1 U2274 ( .A(\REGISTERS[17][28] ), .ZN(n696) );
  INV_X1 U2275 ( .A(\REGISTERS[13][28] ), .ZN(n703) );
  INV_X1 U2276 ( .A(\REGISTERS[9][28] ), .ZN(n706) );
  INV_X1 U2277 ( .A(\REGISTERS[5][28] ), .ZN(n709) );
  INV_X1 U2278 ( .A(\REGISTERS[1][28] ), .ZN(n712) );
  INV_X1 U2279 ( .A(\REGISTERS[29][29] ), .ZN(n653) );
  INV_X1 U2280 ( .A(\REGISTERS[25][29] ), .ZN(n656) );
  INV_X1 U2281 ( .A(\REGISTERS[21][29] ), .ZN(n659) );
  INV_X1 U2282 ( .A(\REGISTERS[17][29] ), .ZN(n662) );
  INV_X1 U2283 ( .A(\REGISTERS[13][29] ), .ZN(n669) );
  INV_X1 U2284 ( .A(\REGISTERS[9][29] ), .ZN(n672) );
  INV_X1 U2285 ( .A(\REGISTERS[5][29] ), .ZN(n675) );
  INV_X1 U2286 ( .A(\REGISTERS[1][29] ), .ZN(n678) );
  INV_X1 U2287 ( .A(\REGISTERS[29][30] ), .ZN(n619) );
  INV_X1 U2288 ( .A(\REGISTERS[25][30] ), .ZN(n622) );
  INV_X1 U2289 ( .A(\REGISTERS[21][30] ), .ZN(n625) );
  INV_X1 U2290 ( .A(\REGISTERS[17][30] ), .ZN(n628) );
  INV_X1 U2291 ( .A(\REGISTERS[13][30] ), .ZN(n635) );
  INV_X1 U2292 ( .A(\REGISTERS[9][30] ), .ZN(n638) );
  INV_X1 U2293 ( .A(\REGISTERS[5][30] ), .ZN(n641) );
  INV_X1 U2294 ( .A(\REGISTERS[1][30] ), .ZN(n644) );
  INV_X1 U2295 ( .A(\REGISTERS[29][31] ), .ZN(n555) );
  INV_X1 U2296 ( .A(\REGISTERS[25][31] ), .ZN(n562) );
  INV_X1 U2297 ( .A(\REGISTERS[21][31] ), .ZN(n569) );
  INV_X1 U2298 ( .A(\REGISTERS[17][31] ), .ZN(n576) );
  INV_X1 U2299 ( .A(\REGISTERS[13][31] ), .ZN(n587) );
  INV_X1 U2300 ( .A(\REGISTERS[9][31] ), .ZN(n594) );
  INV_X1 U2301 ( .A(\REGISTERS[5][31] ), .ZN(n601) );
  INV_X1 U2302 ( .A(\REGISTERS[1][31] ), .ZN(n608) );
  BUF_X1 U2303 ( .A(RESET), .Z(n3094) );
  INV_X1 U2304 ( .A(ADD_RD2[2]), .ZN(n1681) );
  INV_X1 U2305 ( .A(ADD_RD2[1]), .ZN(n1677) );
  INV_X1 U2306 ( .A(ADD_RD1[2]), .ZN(n2305) );
  INV_X1 U2307 ( .A(ADD_RD1[1]), .ZN(n2303) );
  INV_X1 U2308 ( .A(ADD_WR[4]), .ZN(n539) );
  INV_X1 U2309 ( .A(ADD_WR[3]), .ZN(n537) );
endmodule


module D_Reg_generic_N32_10 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net55849, net55850, net55851, net55852, net55853, net55854,
         net55855, net55856, net55857, net55858, net55859, net55860, net55861,
         net55862, net55863, net55864, net55865, net55866, net55867, net55868,
         n48, n33, n34, n35, n36, n37, n38, n42, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n74, n75, n76, n77, n78, n79, n80,
         n81, n82;
  assign n48 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(CLK), .RN(n82), .Q(Q[31]), .QN(net55868)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(CLK), .RN(n80), .Q(Q[30]), .QN(net55867)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(CLK), .RN(n82), .Q(Q[29]), .QN(net55866)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(CLK), .RN(n80), .Q(Q[28]), .QN(net55865)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(CLK), .RN(n82), .Q(Q[27]), .QN(net55864)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(CLK), .RN(n80), .Q(Q[26]), .QN(net55863)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(CLK), .RN(n80), .Q(Q[25]), .QN(net55862)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(CLK), .RN(n80), .Q(Q[24]), .QN(net55861)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(CLK), .RN(n82), .Q(Q[23]), .QN(net55860)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(CLK), .RN(n80), .Q(Q[22]), .QN(net55859)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(CLK), .RN(n80), .Q(Q[21]), .QN(net55858)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(CLK), .RN(n80), .Q(Q[20]), .QN(net55857)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(CLK), .RN(n82), .Q(Q[19]), .QN(net55856)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(CLK), .RN(n81), .Q(Q[18]), .QN(net55855)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(CLK), .RN(n81), .Q(Q[17]), .QN(net55854)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(CLK), .RN(n81), .Q(Q[16]), .QN(net55853)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(CLK), .RN(n80), .Q(Q[15]), .QN(net55852)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(CLK), .RN(n81), .Q(Q[14]), .QN(net55851)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(CLK), .RN(n81), .Q(Q[13]), .QN(net55850)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(CLK), .RN(n81), .Q(Q[12]), .QN(net55849)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(CLK), .RN(n81), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(CLK), .RN(n81), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(CLK), .RN(n82), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(CLK), .RN(n80), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(CLK), .RN(n82), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(CLK), .RN(n80), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(CLK), .RN(n81), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(CLK), .RN(n80), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(CLK), .RN(n81), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(CLK), .RN(n81), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(CLK), .RN(n81), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(CLK), .RN(n82), .Q(Q[0]) );
  BUF_X1 U2 ( .A(n74), .Z(n77) );
  BUF_X1 U3 ( .A(n74), .Z(n76) );
  BUF_X1 U4 ( .A(n75), .Z(n78) );
  BUF_X1 U5 ( .A(n75), .Z(n79) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n74) );
  BUF_X1 U7 ( .A(ENABLE), .Z(n75) );
  OAI21_X1 U8 ( .B1(net55860), .B2(n78), .A(n33), .ZN(n9) );
  NAND2_X1 U9 ( .A1(n79), .A2(D[23]), .ZN(n33) );
  OAI21_X1 U10 ( .B1(net55861), .B2(n77), .A(n34), .ZN(n8) );
  NAND2_X1 U11 ( .A1(D[24]), .A2(n76), .ZN(n34) );
  OAI21_X1 U12 ( .B1(net55862), .B2(n77), .A(n35), .ZN(n7) );
  NAND2_X1 U13 ( .A1(D[25]), .A2(n76), .ZN(n35) );
  OAI21_X1 U14 ( .B1(net55864), .B2(n77), .A(n37), .ZN(n5) );
  NAND2_X1 U15 ( .A1(D[27]), .A2(n76), .ZN(n37) );
  OAI21_X1 U16 ( .B1(net55852), .B2(n78), .A(n57), .ZN(n17) );
  NAND2_X1 U17 ( .A1(D[15]), .A2(n76), .ZN(n57) );
  OAI21_X1 U18 ( .B1(net55856), .B2(n78), .A(n61), .ZN(n13) );
  NAND2_X1 U19 ( .A1(D[19]), .A2(n76), .ZN(n61) );
  OAI21_X1 U20 ( .B1(net55857), .B2(n78), .A(n62), .ZN(n12) );
  NAND2_X1 U21 ( .A1(D[20]), .A2(n76), .ZN(n62) );
  OAI21_X1 U22 ( .B1(net55863), .B2(n78), .A(n36), .ZN(n6) );
  NAND2_X1 U23 ( .A1(D[26]), .A2(n76), .ZN(n36) );
  OAI21_X1 U24 ( .B1(net55865), .B2(n78), .A(n38), .ZN(n4) );
  NAND2_X1 U25 ( .A1(D[28]), .A2(n76), .ZN(n38) );
  OAI21_X1 U26 ( .B1(net55866), .B2(n78), .A(n42), .ZN(n3) );
  NAND2_X1 U27 ( .A1(D[29]), .A2(n76), .ZN(n42) );
  OAI21_X1 U28 ( .B1(net55858), .B2(n79), .A(n63), .ZN(n11) );
  NAND2_X1 U29 ( .A1(D[21]), .A2(n76), .ZN(n63) );
  OAI21_X1 U30 ( .B1(net55859), .B2(n79), .A(n64), .ZN(n10) );
  NAND2_X1 U31 ( .A1(D[22]), .A2(n76), .ZN(n64) );
  OAI21_X1 U32 ( .B1(net55868), .B2(n79), .A(n65), .ZN(n1) );
  NAND2_X1 U33 ( .A1(D[31]), .A2(n76), .ZN(n65) );
  OAI21_X1 U34 ( .B1(net55850), .B2(n77), .A(n55), .ZN(n19) );
  NAND2_X1 U35 ( .A1(D[13]), .A2(n77), .ZN(n55) );
  OAI21_X1 U36 ( .B1(net55867), .B2(n77), .A(n54), .ZN(n2) );
  NAND2_X1 U37 ( .A1(D[30]), .A2(n77), .ZN(n54) );
  OAI21_X1 U38 ( .B1(net55849), .B2(n78), .A(n53), .ZN(n20) );
  NAND2_X1 U39 ( .A1(D[12]), .A2(n77), .ZN(n53) );
  OAI21_X1 U40 ( .B1(net55851), .B2(n78), .A(n56), .ZN(n18) );
  NAND2_X1 U41 ( .A1(D[14]), .A2(n77), .ZN(n56) );
  OAI21_X1 U42 ( .B1(net55853), .B2(n78), .A(n58), .ZN(n16) );
  NAND2_X1 U43 ( .A1(D[16]), .A2(n77), .ZN(n58) );
  OAI21_X1 U44 ( .B1(net55854), .B2(n78), .A(n59), .ZN(n15) );
  NAND2_X1 U45 ( .A1(D[17]), .A2(n77), .ZN(n59) );
  OAI21_X1 U46 ( .B1(net55855), .B2(n78), .A(n60), .ZN(n14) );
  NAND2_X1 U47 ( .A1(D[18]), .A2(n77), .ZN(n60) );
  BUF_X1 U48 ( .A(n48), .Z(n81) );
  BUF_X1 U49 ( .A(n48), .Z(n80) );
  BUF_X1 U50 ( .A(n48), .Z(n82) );
  MUX2_X1 U51 ( .A(Q[0]), .B(D[0]), .S(n79), .Z(n32) );
  MUX2_X1 U52 ( .A(Q[1]), .B(D[1]), .S(n79), .Z(n31) );
  MUX2_X1 U53 ( .A(Q[2]), .B(D[2]), .S(n79), .Z(n30) );
  MUX2_X1 U54 ( .A(Q[3]), .B(D[3]), .S(n79), .Z(n29) );
  MUX2_X1 U55 ( .A(Q[4]), .B(D[4]), .S(n79), .Z(n28) );
  MUX2_X1 U56 ( .A(Q[5]), .B(D[5]), .S(n79), .Z(n27) );
  MUX2_X1 U57 ( .A(Q[6]), .B(D[6]), .S(n79), .Z(n26) );
  MUX2_X1 U58 ( .A(Q[7]), .B(D[7]), .S(n79), .Z(n25) );
  MUX2_X1 U59 ( .A(Q[8]), .B(D[8]), .S(n79), .Z(n24) );
  MUX2_X1 U60 ( .A(Q[9]), .B(D[9]), .S(n79), .Z(n23) );
  MUX2_X1 U61 ( .A(Q[10]), .B(D[10]), .S(n79), .Z(n22) );
  MUX2_X1 U62 ( .A(Q[11]), .B(D[11]), .S(n79), .Z(n21) );
endmodule


module RCA_gen_N12 ( A, B, Ci, S, Co );
  input [11:0] A;
  input [11:0] B;
  output [11:0] S;
  input Ci;
  output Co;

  wire   [11:1] CTMP;

  FA_0 FAI_0 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_523 FAI_1 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_522 FAI_2 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_521 FAI_3 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_520 FAI_4 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_519 FAI_5 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_518 FAI_6 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_517 FAI_7 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_516 FAI_8 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_515 FAI_9 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_514 FAI_10 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_513 FAI_11 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(Co) );
endmodule


module D_Reg_generic_N32_0 ( D, CLK, RESET, ENABLE, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RESET, ENABLE;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, net55767, net55768, net55769, net55770, net55771,
         net55772, net55773, net55774, net55775, net55776, net55777, net55778,
         net55779, net55780, net55781, net55782, net55783, net55784, net55785,
         net55786, net55787, net55788, net55789, net55790, net55791, net55792,
         net55793, net55794, net55795, net55796, net55797, net55798, n41, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n42, n43, n44, n45, n46, n47, n48, n49, n50;
  assign n41 = RESET;

  DFFR_X1 \Q_reg[31]  ( .D(n96), .CK(CLK), .RN(n49), .Q(Q[31]), .QN(net55798)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(CLK), .RN(n49), .Q(Q[30]), .QN(net55797)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(CLK), .RN(n49), .Q(Q[29]), .QN(net55796)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(CLK), .RN(n49), .Q(Q[28]), .QN(net55795)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(CLK), .RN(n49), .Q(Q[27]), .QN(net55794)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(CLK), .RN(n49), .Q(Q[26]), .QN(net55793)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(CLK), .RN(n49), .Q(Q[25]), .QN(net55792)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(CLK), .RN(n49), .Q(Q[24]), .QN(net55791)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(CLK), .RN(n49), .Q(Q[23]), .QN(net55790)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(CLK), .RN(n49), .Q(Q[22]), .QN(net55789)
         );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(CLK), .RN(n49), .Q(Q[21]), .QN(net55788)
         );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(CLK), .RN(n49), .Q(Q[20]), .QN(net55787)
         );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(CLK), .RN(n48), .Q(Q[19]), .QN(net55786)
         );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(CLK), .RN(n48), .Q(Q[18]), .QN(net55785)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(CLK), .RN(n48), .Q(Q[17]), .QN(net55784)
         );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(CLK), .RN(n48), .Q(Q[16]), .QN(net55783)
         );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(CLK), .RN(n48), .Q(Q[15]), .QN(net55782)
         );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(CLK), .RN(n48), .Q(Q[14]), .QN(net55781)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(CLK), .RN(n48), .Q(Q[13]), .QN(net55780)
         );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(CLK), .RN(n48), .Q(Q[12]), .QN(net55779)
         );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(CLK), .RN(n48), .Q(Q[11]), .QN(net55778)
         );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(CLK), .RN(n48), .Q(Q[10]), .QN(net55777)
         );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(CLK), .RN(n48), .Q(Q[9]), .QN(net55776) );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(CLK), .RN(n48), .Q(Q[8]), .QN(net55775) );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(CLK), .RN(n50), .Q(Q[7]), .QN(net55774) );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(CLK), .RN(n50), .Q(Q[6]), .QN(net55773) );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(CLK), .RN(n50), .Q(Q[5]), .QN(net55772) );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(CLK), .RN(n50), .Q(Q[4]), .QN(net55771) );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(CLK), .RN(n50), .Q(Q[3]), .QN(net55770) );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(CLK), .RN(n50), .Q(Q[2]), .QN(net55769) );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(CLK), .RN(n50), .Q(Q[1]), .QN(net55768) );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(CLK), .RN(n50), .Q(Q[0]), .QN(net55767) );
  BUF_X1 U2 ( .A(ENABLE), .Z(n42) );
  BUF_X1 U3 ( .A(ENABLE), .Z(n43) );
  BUF_X1 U4 ( .A(ENABLE), .Z(n44) );
  BUF_X1 U5 ( .A(ENABLE), .Z(n46) );
  BUF_X1 U6 ( .A(ENABLE), .Z(n45) );
  OAI21_X1 U7 ( .B1(net55798), .B2(n45), .A(n1), .ZN(n96) );
  NAND2_X1 U8 ( .A1(n47), .A2(D[31]), .ZN(n1) );
  OAI21_X1 U9 ( .B1(net55768), .B2(n47), .A(n31), .ZN(n66) );
  NAND2_X1 U10 ( .A1(D[1]), .A2(n42), .ZN(n31) );
  OAI21_X1 U11 ( .B1(net55769), .B2(n47), .A(n30), .ZN(n67) );
  NAND2_X1 U12 ( .A1(D[2]), .A2(n42), .ZN(n30) );
  OAI21_X1 U13 ( .B1(net55770), .B2(n47), .A(n29), .ZN(n68) );
  NAND2_X1 U14 ( .A1(D[3]), .A2(n42), .ZN(n29) );
  OAI21_X1 U15 ( .B1(net55791), .B2(n44), .A(n8), .ZN(n89) );
  NAND2_X1 U16 ( .A1(D[24]), .A2(n43), .ZN(n8) );
  OAI21_X1 U17 ( .B1(net55793), .B2(n44), .A(n6), .ZN(n91) );
  NAND2_X1 U18 ( .A1(D[26]), .A2(n43), .ZN(n6) );
  OAI21_X1 U19 ( .B1(net55794), .B2(n44), .A(n5), .ZN(n92) );
  NAND2_X1 U20 ( .A1(D[27]), .A2(n42), .ZN(n5) );
  OAI21_X1 U21 ( .B1(net55796), .B2(n44), .A(n3), .ZN(n94) );
  NAND2_X1 U22 ( .A1(D[29]), .A2(n42), .ZN(n3) );
  OAI21_X1 U23 ( .B1(net55797), .B2(n44), .A(n2), .ZN(n95) );
  NAND2_X1 U24 ( .A1(D[30]), .A2(n42), .ZN(n2) );
  OAI21_X1 U25 ( .B1(net55767), .B2(n45), .A(n32), .ZN(n65) );
  NAND2_X1 U26 ( .A1(D[0]), .A2(n42), .ZN(n32) );
  OAI21_X1 U27 ( .B1(net55771), .B2(n46), .A(n28), .ZN(n69) );
  NAND2_X1 U28 ( .A1(D[4]), .A2(n42), .ZN(n28) );
  OAI21_X1 U29 ( .B1(net55772), .B2(n46), .A(n27), .ZN(n70) );
  NAND2_X1 U30 ( .A1(D[5]), .A2(n42), .ZN(n27) );
  OAI21_X1 U31 ( .B1(net55773), .B2(n46), .A(n26), .ZN(n71) );
  NAND2_X1 U32 ( .A1(D[6]), .A2(n42), .ZN(n26) );
  OAI21_X1 U33 ( .B1(net55774), .B2(n46), .A(n25), .ZN(n72) );
  NAND2_X1 U34 ( .A1(D[7]), .A2(n42), .ZN(n25) );
  OAI21_X1 U35 ( .B1(net55775), .B2(n46), .A(n24), .ZN(n73) );
  NAND2_X1 U36 ( .A1(D[8]), .A2(n43), .ZN(n24) );
  OAI21_X1 U37 ( .B1(net55776), .B2(n46), .A(n23), .ZN(n74) );
  NAND2_X1 U38 ( .A1(D[9]), .A2(n43), .ZN(n23) );
  OAI21_X1 U39 ( .B1(net55777), .B2(n46), .A(n22), .ZN(n75) );
  NAND2_X1 U40 ( .A1(D[10]), .A2(n43), .ZN(n22) );
  OAI21_X1 U41 ( .B1(net55778), .B2(n46), .A(n21), .ZN(n76) );
  NAND2_X1 U42 ( .A1(D[11]), .A2(n43), .ZN(n21) );
  OAI21_X1 U43 ( .B1(net55779), .B2(n46), .A(n20), .ZN(n77) );
  NAND2_X1 U44 ( .A1(D[12]), .A2(n43), .ZN(n20) );
  OAI21_X1 U45 ( .B1(net55780), .B2(n46), .A(n19), .ZN(n78) );
  NAND2_X1 U46 ( .A1(D[13]), .A2(n43), .ZN(n19) );
  OAI21_X1 U47 ( .B1(net55781), .B2(n46), .A(n18), .ZN(n79) );
  NAND2_X1 U48 ( .A1(D[14]), .A2(n43), .ZN(n18) );
  OAI21_X1 U49 ( .B1(net55788), .B2(n45), .A(n11), .ZN(n86) );
  NAND2_X1 U50 ( .A1(D[21]), .A2(n43), .ZN(n11) );
  OAI21_X1 U51 ( .B1(net55790), .B2(n45), .A(n9), .ZN(n88) );
  NAND2_X1 U52 ( .A1(D[23]), .A2(n43), .ZN(n9) );
  OAI21_X1 U53 ( .B1(net55792), .B2(n45), .A(n7), .ZN(n90) );
  NAND2_X1 U54 ( .A1(D[25]), .A2(n43), .ZN(n7) );
  OAI21_X1 U55 ( .B1(net55795), .B2(n45), .A(n4), .ZN(n93) );
  NAND2_X1 U56 ( .A1(D[28]), .A2(n42), .ZN(n4) );
  OAI21_X1 U57 ( .B1(net55782), .B2(n46), .A(n17), .ZN(n80) );
  NAND2_X1 U58 ( .A1(D[15]), .A2(n44), .ZN(n17) );
  OAI21_X1 U59 ( .B1(net55783), .B2(n45), .A(n16), .ZN(n81) );
  NAND2_X1 U60 ( .A1(D[16]), .A2(n44), .ZN(n16) );
  OAI21_X1 U61 ( .B1(net55784), .B2(n45), .A(n15), .ZN(n82) );
  NAND2_X1 U62 ( .A1(D[17]), .A2(n44), .ZN(n15) );
  OAI21_X1 U63 ( .B1(net55785), .B2(n45), .A(n14), .ZN(n83) );
  NAND2_X1 U64 ( .A1(D[18]), .A2(n44), .ZN(n14) );
  OAI21_X1 U65 ( .B1(net55786), .B2(n45), .A(n13), .ZN(n84) );
  NAND2_X1 U66 ( .A1(D[19]), .A2(n44), .ZN(n13) );
  OAI21_X1 U67 ( .B1(net55787), .B2(n45), .A(n12), .ZN(n85) );
  NAND2_X1 U68 ( .A1(D[20]), .A2(n44), .ZN(n12) );
  OAI21_X1 U69 ( .B1(net55789), .B2(n45), .A(n10), .ZN(n87) );
  NAND2_X1 U70 ( .A1(D[22]), .A2(n44), .ZN(n10) );
  BUF_X1 U71 ( .A(n41), .Z(n48) );
  BUF_X1 U72 ( .A(n41), .Z(n49) );
  BUF_X1 U73 ( .A(n41), .Z(n50) );
  CLKBUF_X1 U74 ( .A(ENABLE), .Z(n47) );
endmodule


module D_Reg_generic_N12 ( D, CLK, RESET, ENABLE, Q );
  input [11:0] D;
  output [11:0] Q;
  input CLK, RESET, ENABLE;
  wire   n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n1, n14;
  assign n1 = RESET;

  DFFR_X1 \Q_reg[11]  ( .D(n36), .CK(CLK), .RN(n14), .Q(Q[11]) );
  DFFR_X1 \Q_reg[10]  ( .D(n35), .CK(CLK), .RN(n14), .Q(Q[10]) );
  DFFR_X1 \Q_reg[9]  ( .D(n34), .CK(CLK), .RN(n14), .Q(Q[9]) );
  DFFR_X1 \Q_reg[8]  ( .D(n33), .CK(CLK), .RN(n14), .Q(Q[8]) );
  DFFR_X1 \Q_reg[7]  ( .D(n32), .CK(CLK), .RN(n14), .Q(Q[7]) );
  DFFR_X1 \Q_reg[6]  ( .D(n31), .CK(CLK), .RN(n14), .Q(Q[6]) );
  DFFR_X1 \Q_reg[5]  ( .D(n30), .CK(CLK), .RN(n14), .Q(Q[5]) );
  DFFR_X1 \Q_reg[4]  ( .D(n29), .CK(CLK), .RN(n14), .Q(Q[4]) );
  DFFR_X1 \Q_reg[3]  ( .D(n28), .CK(CLK), .RN(n14), .Q(Q[3]) );
  DFFR_X1 \Q_reg[2]  ( .D(n27), .CK(CLK), .RN(n14), .Q(Q[2]) );
  DFFR_X1 \Q_reg[1]  ( .D(n26), .CK(CLK), .RN(n14), .Q(Q[1]) );
  DFFR_X1 \Q_reg[0]  ( .D(n25), .CK(CLK), .RN(n14), .Q(Q[0]) );
  BUF_X1 U2 ( .A(n1), .Z(n14) );
  MUX2_X1 U3 ( .A(Q[0]), .B(D[0]), .S(ENABLE), .Z(n25) );
  MUX2_X1 U4 ( .A(Q[1]), .B(D[1]), .S(ENABLE), .Z(n26) );
  MUX2_X1 U5 ( .A(Q[2]), .B(D[2]), .S(ENABLE), .Z(n27) );
  MUX2_X1 U6 ( .A(Q[3]), .B(D[3]), .S(ENABLE), .Z(n28) );
  MUX2_X1 U7 ( .A(Q[4]), .B(D[4]), .S(ENABLE), .Z(n29) );
  MUX2_X1 U8 ( .A(Q[5]), .B(D[5]), .S(ENABLE), .Z(n30) );
  MUX2_X1 U9 ( .A(Q[6]), .B(D[6]), .S(ENABLE), .Z(n31) );
  MUX2_X1 U10 ( .A(Q[7]), .B(D[7]), .S(ENABLE), .Z(n32) );
  MUX2_X1 U11 ( .A(Q[8]), .B(D[8]), .S(ENABLE), .Z(n33) );
  MUX2_X1 U12 ( .A(Q[9]), .B(D[9]), .S(ENABLE), .Z(n34) );
  MUX2_X1 U13 ( .A(Q[10]), .B(D[10]), .S(ENABLE), .Z(n35) );
  MUX2_X1 U14 ( .A(Q[11]), .B(D[11]), .S(ENABLE), .Z(n36) );
endmodule


module MUX21_GENERIC_N12_1 ( A, B, S, Y );
  input [11:0] A;
  input [11:0] B;
  output [11:0] Y;
  input S;


  MUX21_931 MUXes_0 ( .A(A[0]), .B(B[0]), .S(S), .Y(Y[0]) );
  MUX21_930 MUXes_1 ( .A(A[1]), .B(B[1]), .S(S), .Y(Y[1]) );
  MUX21_929 MUXes_2 ( .A(A[2]), .B(B[2]), .S(S), .Y(Y[2]) );
  MUX21_928 MUXes_3 ( .A(A[3]), .B(B[3]), .S(S), .Y(Y[3]) );
  MUX21_927 MUXes_4 ( .A(A[4]), .B(B[4]), .S(S), .Y(Y[4]) );
  MUX21_926 MUXes_5 ( .A(A[5]), .B(B[5]), .S(S), .Y(Y[5]) );
  MUX21_925 MUXes_6 ( .A(A[6]), .B(B[6]), .S(S), .Y(Y[6]) );
  MUX21_924 MUXes_7 ( .A(A[7]), .B(B[7]), .S(S), .Y(Y[7]) );
  MUX21_923 MUXes_8 ( .A(A[8]), .B(B[8]), .S(S), .Y(Y[8]) );
  MUX21_922 MUXes_9 ( .A(A[9]), .B(B[9]), .S(S), .Y(Y[9]) );
  MUX21_921 MUXes_10 ( .A(A[10]), .B(B[10]), .S(S), .Y(Y[10]) );
  MUX21_920 MUXes_11 ( .A(A[11]), .B(B[11]), .S(S), .Y(Y[11]) );
endmodule


module MUX21_GENERIC_N12_0 ( A, B, S, Y );
  input [11:0] A;
  input [11:0] B;
  output [11:0] Y;
  input S;
  wire   n1, n2;
  assign n1 = S;

  MUX21_0 MUXes_0 ( .A(A[0]), .B(B[0]), .S(n2), .Y(Y[0]) );
  MUX21_942 MUXes_1 ( .A(A[1]), .B(B[1]), .S(n2), .Y(Y[1]) );
  MUX21_941 MUXes_2 ( .A(A[2]), .B(B[2]), .S(n2), .Y(Y[2]) );
  MUX21_940 MUXes_3 ( .A(A[3]), .B(B[3]), .S(n2), .Y(Y[3]) );
  MUX21_939 MUXes_4 ( .A(A[4]), .B(B[4]), .S(n2), .Y(Y[4]) );
  MUX21_938 MUXes_5 ( .A(A[5]), .B(B[5]), .S(n2), .Y(Y[5]) );
  MUX21_937 MUXes_6 ( .A(A[6]), .B(B[6]), .S(n2), .Y(Y[6]) );
  MUX21_936 MUXes_7 ( .A(A[7]), .B(B[7]), .S(n2), .Y(Y[7]) );
  MUX21_935 MUXes_8 ( .A(A[8]), .B(B[8]), .S(n2), .Y(Y[8]) );
  MUX21_934 MUXes_9 ( .A(A[9]), .B(B[9]), .S(n2), .Y(Y[9]) );
  MUX21_933 MUXes_10 ( .A(A[10]), .B(B[10]), .S(n2), .Y(Y[10]) );
  MUX21_932 MUXes_11 ( .A(A[11]), .B(B[11]), .S(n2), .Y(Y[11]) );
  BUF_X2 U1 ( .A(n1), .Z(n2) );
endmodule


module WritebackUnit_Nbit32 ( WBMux_sel, NPC8, NPC12, DataIn_DMem, DataIn_ALU, 
        WB_DataOut );
  input [1:0] WBMux_sel;
  input [31:0] NPC8;
  input [31:0] NPC12;
  input [31:0] DataIn_DMem;
  input [31:0] DataIn_ALU;
  output [31:0] WB_DataOut;


  mux41_generic_N32_1 WB_MUX ( .A(DataIn_DMem), .B(DataIn_ALU), .C(NPC8), .D(
        NPC12), .S(WBMux_sel), .Y(WB_DataOut) );
endmodule


module MemoryUnit_Nbit32_Addr_bit5 ( CLK, RST, REG_EN_M, DataIn_DMem, 
        DataIn_ALU, DataIn_RegB, WR_Addr_E, DataOut_Load, DataOut_Branch, 
        WB_Address, DataOut_Store, Addr_DMem );
  input [31:0] DataIn_DMem;
  input [31:0] DataIn_ALU;
  input [31:0] DataIn_RegB;
  input [4:0] WR_Addr_E;
  output [31:0] DataOut_Load;
  output [31:0] DataOut_Branch;
  output [4:0] WB_Address;
  output [31:0] DataOut_Store;
  output [9:0] Addr_DMem;
  input CLK, RST, REG_EN_M;
  wire   \DataIn_ALU[9] , \DataIn_ALU[8] , \DataIn_ALU[7] , \DataIn_ALU[6] ,
         \DataIn_ALU[5] , \DataIn_ALU[4] , \DataIn_ALU[3] , \DataIn_ALU[2] ,
         \DataIn_ALU[1] , \DataIn_ALU[0] ;
  assign DataOut_Store[31] = DataIn_RegB[31];
  assign DataOut_Store[30] = DataIn_RegB[30];
  assign DataOut_Store[29] = DataIn_RegB[29];
  assign DataOut_Store[28] = DataIn_RegB[28];
  assign DataOut_Store[27] = DataIn_RegB[27];
  assign DataOut_Store[26] = DataIn_RegB[26];
  assign DataOut_Store[25] = DataIn_RegB[25];
  assign DataOut_Store[24] = DataIn_RegB[24];
  assign DataOut_Store[23] = DataIn_RegB[23];
  assign DataOut_Store[22] = DataIn_RegB[22];
  assign DataOut_Store[21] = DataIn_RegB[21];
  assign DataOut_Store[20] = DataIn_RegB[20];
  assign DataOut_Store[19] = DataIn_RegB[19];
  assign DataOut_Store[18] = DataIn_RegB[18];
  assign DataOut_Store[17] = DataIn_RegB[17];
  assign DataOut_Store[16] = DataIn_RegB[16];
  assign DataOut_Store[15] = DataIn_RegB[15];
  assign DataOut_Store[14] = DataIn_RegB[14];
  assign DataOut_Store[13] = DataIn_RegB[13];
  assign DataOut_Store[12] = DataIn_RegB[12];
  assign DataOut_Store[11] = DataIn_RegB[11];
  assign DataOut_Store[10] = DataIn_RegB[10];
  assign DataOut_Store[9] = DataIn_RegB[9];
  assign DataOut_Store[8] = DataIn_RegB[8];
  assign DataOut_Store[7] = DataIn_RegB[7];
  assign DataOut_Store[6] = DataIn_RegB[6];
  assign DataOut_Store[5] = DataIn_RegB[5];
  assign DataOut_Store[4] = DataIn_RegB[4];
  assign DataOut_Store[3] = DataIn_RegB[3];
  assign DataOut_Store[2] = DataIn_RegB[2];
  assign DataOut_Store[1] = DataIn_RegB[1];
  assign DataOut_Store[0] = DataIn_RegB[0];
  assign Addr_DMem[9] = \DataIn_ALU[9] ;
  assign \DataIn_ALU[9]  = DataIn_ALU[9];
  assign Addr_DMem[8] = \DataIn_ALU[8] ;
  assign \DataIn_ALU[8]  = DataIn_ALU[8];
  assign Addr_DMem[7] = \DataIn_ALU[7] ;
  assign \DataIn_ALU[7]  = DataIn_ALU[7];
  assign Addr_DMem[6] = \DataIn_ALU[6] ;
  assign \DataIn_ALU[6]  = DataIn_ALU[6];
  assign Addr_DMem[5] = \DataIn_ALU[5] ;
  assign \DataIn_ALU[5]  = DataIn_ALU[5];
  assign Addr_DMem[4] = \DataIn_ALU[4] ;
  assign \DataIn_ALU[4]  = DataIn_ALU[4];
  assign Addr_DMem[3] = \DataIn_ALU[3] ;
  assign \DataIn_ALU[3]  = DataIn_ALU[3];
  assign Addr_DMem[2] = \DataIn_ALU[2] ;
  assign \DataIn_ALU[2]  = DataIn_ALU[2];
  assign Addr_DMem[1] = \DataIn_ALU[1] ;
  assign \DataIn_ALU[1]  = DataIn_ALU[1];
  assign Addr_DMem[0] = \DataIn_ALU[0] ;
  assign \DataIn_ALU[0]  = DataIn_ALU[0];

  D_Reg_generic_N32_2 LMD ( .D(DataIn_DMem), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_M), .Q(DataOut_Load) );
  D_Reg_generic_N32_1 BRANCH_REG ( .D({DataIn_ALU[31:10], \DataIn_ALU[9] , 
        \DataIn_ALU[8] , \DataIn_ALU[7] , \DataIn_ALU[6] , \DataIn_ALU[5] , 
        \DataIn_ALU[4] , \DataIn_ALU[3] , \DataIn_ALU[2] , \DataIn_ALU[1] , 
        \DataIn_ALU[0] }), .CLK(CLK), .RESET(RST), .ENABLE(REG_EN_M), .Q(
        DataOut_Branch) );
  D_Reg_generic_N5_1 REGWR ( .D(WR_Addr_E), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_M), .Q(WB_Address) );
endmodule


module ExecutionUnit_Nbit32_Addr_bit5 ( CLK, RST, REG_EN_E, MuxA_Sel, MuxB_Sel, 
        ALU_Config, Sign, BrCond, AddrComp, NPC_In, DataA, DataB, DataIMM, 
        Wr_Addr_D, NPC_Out, ALU_Out, DataBtoDMem, J_addr, Wr_Addr_E, Br_taken
 );
  input [1:0] MuxA_Sel;
  input [1:0] MuxB_Sel;
  input [4:0] ALU_Config;
  input [1:0] BrCond;
  input [31:0] NPC_In;
  input [31:0] DataA;
  input [31:0] DataB;
  input [31:0] DataIMM;
  input [4:0] Wr_Addr_D;
  output [31:0] NPC_Out;
  output [31:0] ALU_Out;
  output [31:0] DataBtoDMem;
  output [31:0] J_addr;
  output [4:0] Wr_Addr_E;
  input CLK, RST, REG_EN_E, Sign, AddrComp;
  output Br_taken;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [31:0] Op1;
  wire   [31:0] Op2;
  assign n2 = DataB[2];
  assign n3 = DataB[1];
  assign n4 = NPC_In[2];
  assign n5 = DataB[0];
  assign n6 = DataA[1];
  assign n7 = NPC_In[1];

  Br_Comp_Nbit32 BrZ ( .A({DataA[31:2], n12, DataA[0]}), .Br_cond(BrCond), 
        .Taken(Br_taken) );
  mux41_generic_N32_3 MUXA ( .A({NPC_In[31:3], n4, n7, NPC_In[0]}), .B({
        DataA[31:2], n6, DataA[0]}), .C({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .D({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .S(MuxA_Sel), .Y({Op1[31:18], n10, Op1[16], n1, Op1[14:8], n9, n8, 
        Op1[5:0]}) );
  mux41_generic_N32_2 MUXB ( .A({DataB[31:3], n2, n3, n5}), .B(DataIMM), .C({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .S(MuxB_Sel), .Y(Op2) );
  ALU_N32 ALUnit ( .FUNC(ALU_Config), .Sign(Sign), .AddrComp(AddrComp), 
        .DATA1({Op1[31:18], n10, Op1[16], n1, Op1[14:11], n17, Op1[9:8], n9, 
        n8, Op1[5:0]}), .DATA2(Op2), .OUTALU(J_addr) );
  D_Reg_generic_N32_5 REGNPC ( .D({NPC_In[31:7], n11, NPC_In[5:3], n4, n13, 
        NPC_In[0]}), .CLK(CLK), .RESET(RST), .ENABLE(REG_EN_E), .Q(NPC_Out) );
  D_Reg_generic_N32_4 REGALU ( .D(J_addr), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_E), .Q(ALU_Out) );
  D_Reg_generic_N32_3 REGB ( .D({DataB[31:4], n15, n14, n16, n5}), .CLK(CLK), 
        .RESET(RST), .ENABLE(REG_EN_E), .Q(DataBtoDMem) );
  D_Reg_generic_N5_2 REGWR ( .D(Wr_Addr_D), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_E), .Q(Wr_Addr_E) );
  CLKBUF_X1 U3 ( .A(NPC_In[6]), .Z(n11) );
  CLKBUF_X1 U4 ( .A(n6), .Z(n12) );
  CLKBUF_X1 U5 ( .A(n7), .Z(n13) );
  CLKBUF_X1 U6 ( .A(n2), .Z(n14) );
  CLKBUF_X1 U7 ( .A(DataB[3]), .Z(n15) );
  CLKBUF_X1 U8 ( .A(n3), .Z(n16) );
  BUF_X2 U9 ( .A(Op1[10]), .Z(n17) );
endmodule


module DecodeUnit_Nbit32_Addr_bit5 ( CLK, RST, RF_RD1, RF_RD2, RF_WR, REG_EN_D, 
        MuxIMM_Sel, MuxRd_Sel, InstrToDecode, NPCin, WB_Data, WB_Addr, DataA, 
        DataB, DataIMM, NPCout, Jr_addr, Wr_Addr_D );
  input [1:0] MuxIMM_Sel;
  input [1:0] MuxRd_Sel;
  input [31:0] InstrToDecode;
  input [31:0] NPCin;
  input [31:0] WB_Data;
  input [4:0] WB_Addr;
  output [31:0] DataA;
  output [31:0] DataB;
  output [31:0] DataIMM;
  output [31:0] NPCout;
  output [31:0] Jr_addr;
  output [4:0] Wr_Addr_D;
  input CLK, RST, RF_RD1, RF_RD2, RF_WR, REG_EN_D;
  wire   RF_EN;
  wire   [31:0] RF_outB;
  wire   [4:0] WRaddr;
  wire   [31:0] MuxIMM_Out;

  register_file_gen_Nbit32_Nreg32 REG_FILE ( .RESET(RST), .ENABLE(RF_EN), .WR(
        RF_WR), .RD1(RF_RD1), .RD2(RF_RD2), .ADD_WR(WB_Addr), .ADD_RD1(
        InstrToDecode[25:21]), .ADD_RD2(InstrToDecode[20:16]), .DATAIN(WB_Data), .OUT1(Jr_addr), .OUT2(RF_outB) );
  mux41_generic_N5 MUXWR ( .A(InstrToDecode[20:16]), .B(InstrToDecode[15:11]), 
        .C({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .S(MuxRd_Sel), .Y(WRaddr) );
  mux41_generic_N32_0 MUXIMM ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        InstrToDecode[15:0]}), .B({InstrToDecode[15], InstrToDecode[15], 
        InstrToDecode[15], InstrToDecode[15], InstrToDecode[15], 
        InstrToDecode[15], InstrToDecode[15], InstrToDecode[15], 
        InstrToDecode[15], InstrToDecode[15], InstrToDecode[15], 
        InstrToDecode[15], InstrToDecode[15], InstrToDecode[15], 
        InstrToDecode[15], InstrToDecode[15], InstrToDecode[15:0]}), .C({
        InstrToDecode[15:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({
        InstrToDecode[25], InstrToDecode[25], InstrToDecode[25], 
        InstrToDecode[25], InstrToDecode[25], InstrToDecode[25], 
        InstrToDecode[25:0]}), .S(MuxIMM_Sel), .Y(MuxIMM_Out) );
  D_Reg_generic_N32_9 REGA ( .D(Jr_addr), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_D), .Q(DataA) );
  D_Reg_generic_N32_8 REGB ( .D(RF_outB), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_D), .Q(DataB) );
  D_Reg_generic_N32_7 REGIMM ( .D(MuxIMM_Out), .CLK(CLK), .RESET(RST), 
        .ENABLE(REG_EN_D), .Q(DataIMM) );
  D_Reg_generic_N32_6 REGNPC ( .D(NPCin), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_D), .Q(NPCout) );
  D_Reg_generic_N5_0 REGWR ( .D(WRaddr), .CLK(CLK), .RESET(RST), .ENABLE(
        REG_EN_D), .Q(Wr_Addr_D) );
  OR2_X1 U3 ( .A1(REG_EN_D), .A2(RF_WR), .ZN(RF_EN) );
endmodule


module FetchUnit_Nbit32_Iram_bit12 ( CLK, RST, IR_EN, NPC_EN, PC_EN, Jr_Sel, 
        J_Sel, Br_taken, Jr_addr, J_addr, IMem_Instr, InstrToDecode, 
        NPCToDecode, IMem_Addr, Opcode, Func );
  input [11:0] Jr_addr;
  input [11:0] J_addr;
  input [31:0] IMem_Instr;
  output [31:0] InstrToDecode;
  output [31:0] NPCToDecode;
  output [11:0] IMem_Addr;
  output [5:0] Opcode;
  output [10:0] Func;
  input CLK, RST, IR_EN, NPC_EN, PC_EN, Jr_Sel, J_Sel, Br_taken;
  wire   \IMem_Instr[31] , \IMem_Instr[30] , \IMem_Instr[29] ,
         \IMem_Instr[28] , \IMem_Instr[27] , \IMem_Instr[26] ,
         \IMem_Instr[10] , \IMem_Instr[9] , \IMem_Instr[8] , \IMem_Instr[7] ,
         \IMem_Instr[6] , \IMem_Instr[5] , \IMem_Instr[4] , \IMem_Instr[3] ,
         \IMem_Instr[2] , \IMem_Instr[1] , \IMem_Instr[0] , J_Br_Sel;
  wire   [11:0] NPC_input;
  wire   [11:0] JRtoJ_PC;
  wire   [11:0] JtoPC;
  assign Opcode[5] = \IMem_Instr[31] ;
  assign \IMem_Instr[31]  = IMem_Instr[31];
  assign Opcode[4] = \IMem_Instr[30] ;
  assign \IMem_Instr[30]  = IMem_Instr[30];
  assign Opcode[3] = \IMem_Instr[29] ;
  assign \IMem_Instr[29]  = IMem_Instr[29];
  assign Opcode[2] = \IMem_Instr[28] ;
  assign \IMem_Instr[28]  = IMem_Instr[28];
  assign Opcode[1] = \IMem_Instr[27] ;
  assign \IMem_Instr[27]  = IMem_Instr[27];
  assign Opcode[0] = \IMem_Instr[26] ;
  assign \IMem_Instr[26]  = IMem_Instr[26];
  assign Func[10] = \IMem_Instr[10] ;
  assign \IMem_Instr[10]  = IMem_Instr[10];
  assign Func[9] = \IMem_Instr[9] ;
  assign \IMem_Instr[9]  = IMem_Instr[9];
  assign Func[8] = \IMem_Instr[8] ;
  assign \IMem_Instr[8]  = IMem_Instr[8];
  assign Func[7] = \IMem_Instr[7] ;
  assign \IMem_Instr[7]  = IMem_Instr[7];
  assign Func[6] = \IMem_Instr[6] ;
  assign \IMem_Instr[6]  = IMem_Instr[6];
  assign Func[5] = \IMem_Instr[5] ;
  assign \IMem_Instr[5]  = IMem_Instr[5];
  assign Func[4] = \IMem_Instr[4] ;
  assign \IMem_Instr[4]  = IMem_Instr[4];
  assign Func[3] = \IMem_Instr[3] ;
  assign \IMem_Instr[3]  = IMem_Instr[3];
  assign Func[2] = \IMem_Instr[2] ;
  assign \IMem_Instr[2]  = IMem_Instr[2];
  assign Func[1] = \IMem_Instr[1] ;
  assign \IMem_Instr[1]  = IMem_Instr[1];
  assign Func[0] = \IMem_Instr[0] ;
  assign \IMem_Instr[0]  = IMem_Instr[0];

  MUX21_GENERIC_N12_0 MuxJR ( .A(NPC_input), .B(Jr_addr), .S(Jr_Sel), .Y(
        JRtoJ_PC) );
  MUX21_GENERIC_N12_1 MuxJ ( .A(JRtoJ_PC), .B(J_addr), .S(J_Br_Sel), .Y(JtoPC)
         );
  D_Reg_generic_N12 PC ( .D(JtoPC), .CLK(CLK), .RESET(RST), .ENABLE(PC_EN), 
        .Q(IMem_Addr) );
  D_Reg_generic_N32_0 IR ( .D({\IMem_Instr[31] , \IMem_Instr[30] , 
        \IMem_Instr[29] , \IMem_Instr[28] , \IMem_Instr[27] , \IMem_Instr[26] , 
        IMem_Instr[25:11], \IMem_Instr[10] , \IMem_Instr[9] , \IMem_Instr[8] , 
        \IMem_Instr[7] , \IMem_Instr[6] , \IMem_Instr[5] , \IMem_Instr[4] , 
        \IMem_Instr[3] , \IMem_Instr[2] , \IMem_Instr[1] , \IMem_Instr[0] }), 
        .CLK(CLK), .RESET(RST), .ENABLE(IR_EN), .Q(InstrToDecode) );
  RCA_gen_N12 ADDER ( .A(IMem_Addr), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .Ci(1'b0), .S(NPC_input) );
  D_Reg_generic_N32_10 NPC ( .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, NPC_input}), .CLK(CLK), .RESET(RST), .ENABLE(NPC_EN), .Q(
        NPCToDecode) );
  OR2_X1 U3 ( .A1(Br_taken), .A2(J_Sel), .ZN(J_Br_Sel) );
endmodule


module Datapath ( CLK, RST, Opcode, Func, F_PC_EN, F_NPC_EN, F_IR_EN, F_Jr_Sel, 
        F_J_Sel, IMem_Instr, IMem_Addr, D_REG_EN, D_RF_RD1, D_RF_RD2, D_RF_WR, 
        D_IMM_Sel, D_Rd_Sel, E_REG_EN, E_MuxA_Sel, E_MuxB_Sel, E_ALU_Conf, 
        E_Signed, E_BrCond, E_AddrComp, M_REG_EN, DMem_DataOut, DMem_DataIn, 
        DMem_Addr, WB_Mux_sel );
  output [5:0] Opcode;
  output [10:0] Func;
  input [31:0] IMem_Instr;
  output [11:0] IMem_Addr;
  input [1:0] D_IMM_Sel;
  input [1:0] D_Rd_Sel;
  input [1:0] E_MuxA_Sel;
  input [1:0] E_MuxB_Sel;
  input [4:0] E_ALU_Conf;
  input [1:0] E_BrCond;
  input [31:0] DMem_DataOut;
  output [31:0] DMem_DataIn;
  output [9:0] DMem_Addr;
  input [1:0] WB_Mux_sel;
  input CLK, RST, F_PC_EN, F_NPC_EN, F_IR_EN, F_Jr_Sel, F_J_Sel, D_REG_EN,
         D_RF_RD1, D_RF_RD2, D_RF_WR, E_REG_EN, E_Signed, E_AddrComp, M_REG_EN;
  wire   EtoF_Br_taken, n1, n2, n3, n4, n5, n6;
  wire   [31:0] FtoD_instr;
  wire   [31:0] FtoD_NPC;
  wire   [11:0] EtoF_Jaddr;
  wire   [11:0] DtoF_Jraddr;
  wire   [31:0] WtoD_WRdata;
  wire   [4:0] MtoD_WRaddr;
  wire   [31:0] DtoE_DataA;
  wire   [31:0] DtoE_DataB;
  wire   [31:0] DtoE_imm;
  wire   [31:0] DtoE_NPC;
  wire   [4:0] DtoE_WRaddr;
  wire   [31:0] EtoW_NPC;
  wire   [31:0] EtoM_DataALU;
  wire   [31:0] EtoM_DataB;
  wire   [4:0] EtoM_WRaddr;
  wire   [31:0] MtoW_DataMem;
  wire   [31:0] MtoW_DataALU;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39;

  FetchUnit_Nbit32_Iram_bit12 FU ( .CLK(CLK), .RST(RST), .IR_EN(F_IR_EN), 
        .NPC_EN(F_NPC_EN), .PC_EN(F_PC_EN), .Jr_Sel(F_Jr_Sel), .J_Sel(F_J_Sel), 
        .Br_taken(EtoF_Br_taken), .Jr_addr(DtoF_Jraddr), .J_addr(EtoF_Jaddr), 
        .IMem_Instr(IMem_Instr), .InstrToDecode(FtoD_instr), .NPCToDecode(
        FtoD_NPC), .IMem_Addr(IMem_Addr), .Opcode(Opcode), .Func(Func) );
  DecodeUnit_Nbit32_Addr_bit5 DU ( .CLK(CLK), .RST(RST), .RF_RD1(D_RF_RD1), 
        .RF_RD2(D_RF_RD2), .RF_WR(D_RF_WR), .REG_EN_D(D_REG_EN), .MuxIMM_Sel(
        D_IMM_Sel), .MuxRd_Sel(D_Rd_Sel), .InstrToDecode(FtoD_instr), .NPCin(
        FtoD_NPC), .WB_Data(WtoD_WRdata), .WB_Addr(MtoD_WRaddr), .DataA(
        DtoE_DataA), .DataB(DtoE_DataB), .DataIMM(DtoE_imm), .NPCout({
        DtoE_NPC[31:5], n3, n2, DtoE_NPC[2], n4, n1}), .Jr_addr({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, DtoF_Jraddr}), 
        .Wr_Addr_D(DtoE_WRaddr) );
  ExecutionUnit_Nbit32_Addr_bit5 EXU ( .CLK(CLK), .RST(RST), .REG_EN_E(
        E_REG_EN), .MuxA_Sel(E_MuxA_Sel), .MuxB_Sel(E_MuxB_Sel), .ALU_Config(
        E_ALU_Conf), .Sign(E_Signed), .BrCond(E_BrCond), .AddrComp(E_AddrComp), 
        .NPC_In({DtoE_NPC[31:5], n3, n2, DtoE_NPC[2], n4, n1}), .DataA(
        DtoE_DataA), .DataB(DtoE_DataB), .DataIMM(DtoE_imm), .Wr_Addr_D(
        DtoE_WRaddr), .NPC_Out(EtoW_NPC), .ALU_Out(EtoM_DataALU), 
        .DataBtoDMem(EtoM_DataB), .J_addr({SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, EtoF_Jaddr}), .Wr_Addr_E(EtoM_WRaddr), 
        .Br_taken(EtoF_Br_taken) );
  MemoryUnit_Nbit32_Addr_bit5 MEMU ( .CLK(CLK), .RST(RST), .REG_EN_M(M_REG_EN), 
        .DataIn_DMem(DMem_DataOut), .DataIn_ALU(EtoM_DataALU), .DataIn_RegB(
        EtoM_DataB), .WR_Addr_E(EtoM_WRaddr), .DataOut_Load(MtoW_DataMem), 
        .DataOut_Branch(MtoW_DataALU), .WB_Address(MtoD_WRaddr), 
        .DataOut_Store(DMem_DataIn), .Addr_DMem(DMem_Addr) );
  WritebackUnit_Nbit32 WBU ( .WBMux_sel(WB_Mux_sel), .NPC8(EtoW_NPC), .NPC12({
        DtoE_NPC[31:9], n6, DtoE_NPC[7:5], n3, n2, DtoE_NPC[2], n5, n1}), 
        .DataIn_DMem(MtoW_DataMem), .DataIn_ALU(MtoW_DataALU), .WB_DataOut(
        WtoD_WRdata) );
  CLKBUF_X1 U1 ( .A(n4), .Z(n5) );
  CLKBUF_X1 U2 ( .A(DtoE_NPC[8]), .Z(n6) );
endmodule

